magic
tech sky130A
magscale 1 2
timestamp 1725793971
<< dnwell >>
rect 9664 4112 28180 6613
rect 4523 -10546 28180 4112
<< nwell >>
rect 9584 6407 28290 6723
rect 9584 4221 9870 6407
rect 4413 3905 9870 4221
rect 4413 -10340 4729 3905
rect 5580 -6850 7048 -6593
rect 4952 -6902 5590 -6850
rect 5422 -10340 6464 -10054
rect 27974 -10340 28290 6407
rect 4413 -10656 28290 -10340
<< psubdiff >>
rect 4253 6865 4313 6899
rect 28379 6865 28439 6899
rect 4253 6839 4287 6865
rect 28405 6839 28439 6865
rect 4253 -10741 4287 -10715
rect 28405 -10741 28439 -10715
rect 4253 -10775 4313 -10741
rect 28379 -10775 28439 -10741
<< mvnsubdiff >>
rect 9650 6636 28223 6656
rect 9650 6602 9715 6636
rect 28143 6602 28223 6636
rect 9650 6582 28223 6602
rect 9650 6564 9724 6582
rect 9650 4170 9671 6564
rect 9705 4170 9724 6564
rect 9650 4155 9724 4170
rect 4480 4135 9724 4155
rect 4480 4101 4560 4135
rect 9621 4101 9724 4135
rect 4480 4081 9724 4101
rect 28149 6576 28223 6582
rect 4480 4057 4554 4081
rect 4480 -10482 4500 4057
rect 4534 -10482 4554 4057
rect 4480 -10515 4554 -10482
rect 28149 -10509 28169 6576
rect 28203 -10509 28223 6576
rect 28149 -10515 28223 -10509
rect 4480 -10535 28223 -10515
rect 4480 -10569 4560 -10535
rect 28143 -10569 28223 -10535
rect 4480 -10589 28223 -10569
<< psubdiffcont >>
rect 4313 6865 28379 6899
rect 4253 -10715 4287 6839
rect 28405 -10715 28439 6839
rect 4313 -10775 28379 -10741
<< mvnsubdiffcont >>
rect 9715 6602 28143 6636
rect 9671 4170 9705 6564
rect 4560 4101 9621 4135
rect 4500 -10482 4534 4057
rect 28169 -10509 28203 6576
rect 4560 -10569 28143 -10535
<< locali >>
rect 4253 6865 4313 6899
rect 28379 6865 28439 6899
rect 4253 6839 4427 6865
rect 4287 6817 4427 6839
rect 28261 6839 28439 6865
rect 28261 6817 28405 6839
rect 4287 6786 28405 6817
rect 4287 6767 4356 6786
rect 4320 -10614 4356 6767
rect 6872 6292 7410 6786
rect 28327 6778 28405 6786
rect 9650 6644 28223 6656
rect 9650 6594 9678 6644
rect 28150 6594 28223 6644
rect 9650 6579 28223 6594
rect 9671 6564 9705 6579
rect 6087 5973 6255 5990
rect 6087 5872 6108 5973
rect 6233 5872 6255 5973
rect 6087 5856 6255 5872
rect 8199 5973 8367 5990
rect 8199 5872 8220 5973
rect 8345 5872 8367 5973
rect 8199 5856 8367 5872
rect 4466 5261 4537 5274
rect 4466 4869 4475 5261
rect 4528 4869 4537 5261
rect 4466 4856 4537 4869
rect 6576 5266 6647 5280
rect 6576 4876 6587 5266
rect 6636 4876 6647 5266
rect 6576 4862 6647 4876
rect 28149 6576 28223 6579
rect 28149 6530 28169 6576
rect 28203 6530 28223 6576
rect 4481 4143 9617 4159
rect 4481 4135 4582 4143
rect 9580 4135 9617 4143
rect 9671 4135 9705 4170
rect 4481 4126 4560 4135
rect 4481 -10527 4496 4126
rect 4539 4101 4560 4126
rect 9621 4101 9705 4135
rect 9869 6395 27203 6406
rect 9869 6358 27229 6395
rect 4539 4098 4582 4101
rect 9580 4098 9617 4101
rect 4539 4075 9617 4098
rect 4539 -6694 4552 4075
rect 4888 3834 8199 3959
rect 9869 3879 9893 6358
rect 4888 715 5013 3834
rect 5119 3474 5551 3710
rect 5119 3142 5551 3378
rect 7519 3308 7951 3545
rect 5119 2810 5551 3046
rect 7519 2976 7951 3213
rect 5119 2478 5551 2714
rect 7519 2644 7951 2881
rect 5119 2146 5551 2382
rect 7519 2312 7951 2549
rect 5119 1814 5551 2050
rect 7519 1980 7951 2217
rect 5119 1482 5551 1718
rect 7519 1648 7951 1885
rect 5119 1150 5551 1386
rect 7519 1316 7951 1553
rect 5119 818 5551 1054
rect 7519 984 7951 1221
rect 7519 818 7951 889
rect 8074 715 8199 3834
rect 4888 522 8199 715
rect 4888 -5561 5013 522
rect 5117 181 5549 417
rect 5117 -151 5549 85
rect 7517 15 7949 252
rect 5117 -483 5549 -247
rect 7517 -317 7949 -80
rect 5117 -815 5549 -579
rect 7517 -649 7949 -412
rect 5117 -1147 5549 -911
rect 7517 -981 7949 -744
rect 5117 -1479 5549 -1243
rect 7517 -1313 7949 -1076
rect 5117 -1811 5549 -1575
rect 7517 -1645 7949 -1408
rect 5117 -2143 5549 -1907
rect 7517 -1977 7949 -1740
rect 5117 -2475 5549 -2239
rect 7517 -2309 7949 -2072
rect 5117 -2807 5549 -2571
rect 7517 -2641 7949 -2404
rect 5117 -3139 5549 -2903
rect 7517 -2973 7949 -2736
rect 5117 -3471 5549 -3235
rect 7517 -3305 7949 -3068
rect 5117 -3803 5549 -3567
rect 7517 -3637 7949 -3400
rect 5117 -4135 5549 -3899
rect 7517 -3969 7949 -3732
rect 5117 -4467 5549 -4231
rect 7517 -4301 7949 -4064
rect 5117 -4799 5549 -4563
rect 7517 -4633 7949 -4396
rect 5117 -5131 5549 -4895
rect 7517 -4965 7949 -4728
rect 5117 -5463 5549 -5227
rect 7517 -5297 7949 -5060
rect 7517 -5462 7949 -5392
rect 8074 -5560 8199 522
rect 5047 -5561 8199 -5560
rect 4854 -5607 8199 -5561
rect 4854 -5673 5080 -5607
rect 7920 -5673 8199 -5607
rect 4854 -5687 8199 -5673
rect 4854 -5954 5063 -5687
rect 5555 -5798 7091 -5782
rect 5555 -5863 7092 -5798
rect 5555 -5900 5653 -5863
rect 4855 -5976 5062 -5954
rect 4855 -6488 4873 -5976
rect 5044 -6488 5062 -5976
rect 4855 -6504 5062 -6488
rect 5556 -6602 5653 -5900
rect 5702 -5865 7092 -5863
rect 5702 -5900 6076 -5865
rect 5702 -6495 5724 -5900
rect 6049 -6495 6076 -5900
rect 5702 -6602 6076 -6495
rect 6125 -5870 7092 -5865
rect 6125 -5900 6504 -5870
rect 6125 -6495 6145 -5900
rect 6479 -6495 6504 -5900
rect 6125 -6602 6504 -6495
rect 6553 -5900 7092 -5870
rect 6553 -6495 6575 -5900
rect 6954 -6495 7092 -5900
rect 9870 -5966 9893 3879
rect 9866 -6002 9893 -5966
rect 9956 6262 13341 6358
rect 9956 -5966 9989 6262
rect 13318 -5966 13341 6262
rect 9956 -6002 13341 -5966
rect 13404 6262 16789 6358
rect 13404 -5966 13437 6262
rect 16766 -5966 16789 6262
rect 13404 -6002 16789 -5966
rect 16852 6262 20237 6358
rect 16852 -5966 16885 6262
rect 20214 -5966 20237 6262
rect 16852 -6002 20237 -5966
rect 20300 6262 23685 6358
rect 20300 -5966 20333 6262
rect 23662 -5966 23685 6262
rect 20300 -6002 23685 -5966
rect 23748 6262 27133 6358
rect 23748 -5966 23781 6262
rect 27110 -5966 27133 6262
rect 23748 -6002 27133 -5966
rect 27196 -6002 27229 6358
rect 9866 -6035 27229 -6002
rect 9866 -6110 27141 -6035
rect 6553 -6602 7092 -6495
rect 28149 -6188 28162 6530
rect 28207 -6188 28223 6530
rect 28149 -6536 28169 -6188
rect 5556 -6694 7092 -6602
rect 4539 -6783 21805 -6694
rect 4539 -6879 4763 -6783
rect 21770 -6879 21805 -6783
rect 4539 -6934 21805 -6879
rect 22058 -6782 27804 -6698
rect 22058 -6878 22082 -6782
rect 27742 -6878 27804 -6782
rect 4539 -6953 12927 -6934
rect 4539 -10527 4552 -6953
rect 4789 -7552 4903 -6953
rect 6932 -7556 7060 -6953
rect 9081 -7533 9208 -6953
rect 11223 -7558 11360 -6953
rect 12952 -7549 13087 -6934
rect 15286 -7550 15412 -6934
rect 17440 -7556 17566 -6934
rect 19584 -7548 19716 -6934
rect 22058 -6941 27804 -6878
rect 22058 -7051 26600 -6941
rect 26958 -6948 27804 -6941
rect 26958 -7004 27356 -6948
rect 27378 -6952 27804 -6948
rect 26958 -7051 27354 -7004
rect 22058 -7086 27354 -7051
rect 22164 -7435 22595 -7200
rect 27100 -7562 27354 -7086
rect 4776 -7843 4917 -7841
rect 4776 -7994 4919 -7843
rect 4776 -9961 4809 -7994
rect 4857 -8823 4919 -7994
rect 6917 -8628 7239 -7831
rect 8123 -7848 8414 -7832
rect 8123 -7988 8557 -7848
rect 8123 -8628 8454 -7988
rect 6917 -8823 8454 -8628
rect 4857 -8887 8454 -8823
rect 4857 -9961 4917 -8887
rect 6906 -8888 8454 -8887
rect 5382 -9014 6446 -8989
rect 5382 -9932 5410 -9014
rect 4776 -10082 4917 -9961
rect 5381 -9992 5410 -9932
rect 5454 -9071 6446 -9014
rect 5454 -9942 5533 -9071
rect 5574 -9747 5645 -9071
rect 5997 -9754 6068 -9071
rect 6352 -9942 6446 -9071
rect 5454 -9992 6446 -9942
rect 5381 -10017 6446 -9992
rect 5383 -10018 6446 -10017
rect 6906 -9474 7239 -8888
rect 6906 -10049 7233 -9474
rect 8117 -9475 8454 -8888
rect 7544 -10049 7598 -9657
rect 7985 -10049 8039 -9657
rect 8119 -9958 8454 -9475
rect 8497 -9020 8557 -7988
rect 10155 -7989 10427 -7791
rect 10155 -7991 10333 -7989
rect 10155 -9020 10217 -7991
rect 8497 -9136 10217 -9020
rect 8497 -9188 8577 -9136
rect 9616 -9188 10217 -9136
rect 8497 -9311 10217 -9188
rect 8497 -9897 8766 -9311
rect 9132 -9897 9217 -9311
rect 9576 -9897 9661 -9311
rect 10031 -9897 10217 -9311
rect 8497 -9958 10217 -9897
rect 8119 -9961 10217 -9958
rect 10260 -9961 10333 -7991
rect 10376 -9016 10427 -7989
rect 12764 -7842 12894 -7816
rect 12764 -7985 13018 -7842
rect 12764 -7989 12929 -7985
rect 10376 -9019 10480 -9016
rect 10376 -9589 10557 -9019
rect 12764 -9589 12813 -7989
rect 10376 -9773 12813 -9589
rect 10376 -9961 10557 -9773
rect 8119 -10049 10557 -9961
rect 6906 -10082 10557 -10049
rect 12764 -9978 12813 -9773
rect 12856 -9963 12929 -7989
rect 12972 -9963 13018 -7985
rect 12856 -9978 13018 -9963
rect 12764 -10082 13018 -9978
rect 15034 -7987 15164 -7848
rect 15034 -9978 15077 -7987
rect 15120 -9978 15164 -7987
rect 15034 -10082 15164 -9978
rect 17131 -7983 17217 -7834
rect 17131 -9958 17151 -7983
rect 17194 -9958 17217 -7983
rect 17131 -10082 17217 -9958
rect 19277 -7985 19363 -7841
rect 19277 -9955 19295 -7985
rect 19338 -9955 19363 -7985
rect 19277 -10082 19363 -9955
rect 21426 -7985 21512 -7841
rect 21426 -9949 21449 -7985
rect 21492 -9949 21512 -7985
rect 21426 -10082 21512 -9949
rect 23572 -7985 23658 -7836
rect 23572 -9949 23593 -7985
rect 23636 -9949 23658 -7985
rect 23572 -10082 23658 -9949
rect 25772 -7987 25896 -7838
rect 25772 -9966 25808 -7987
rect 25851 -9966 25896 -7987
rect 25772 -10082 25896 -9966
rect 4690 -10161 27989 -10082
rect 4690 -10256 4763 -10161
rect 27915 -10256 27989 -10161
rect 4690 -10389 27989 -10256
rect 4690 -10488 5783 -10389
rect 4481 -10530 4552 -10527
rect 28203 -6536 28223 -6188
rect 28169 -10530 28203 -10509
rect 4481 -10535 28227 -10530
rect 4481 -10569 4560 -10535
rect 28143 -10550 28227 -10535
rect 4481 -10595 4595 -10569
rect 28200 -10595 28227 -10550
rect 4481 -10613 28227 -10595
rect 4287 -10665 4356 -10614
rect 28327 -10618 28361 6778
rect 28327 -10665 28405 -10618
rect 4287 -10704 28405 -10665
rect 4287 -10715 4386 -10704
rect 4253 -10741 4386 -10715
rect 28323 -10715 28405 -10704
rect 28323 -10741 28439 -10715
rect 4253 -10775 4313 -10741
rect 28379 -10775 28439 -10741
<< viali >>
rect 4427 6865 28261 6871
rect 4427 6817 28261 6865
rect 4270 -10614 4287 6767
rect 4287 -10614 4320 6767
rect 9678 6636 28150 6644
rect 9678 6602 9715 6636
rect 9715 6602 28143 6636
rect 28143 6602 28150 6636
rect 9678 6594 28150 6602
rect 6108 5872 6233 5973
rect 8220 5872 8345 5973
rect 4475 4869 4528 5261
rect 6587 4876 6636 5266
rect 4582 4135 9580 4143
rect 4496 4057 4539 4126
rect 4582 4101 9580 4135
rect 4582 4098 9580 4101
rect 4496 -10482 4500 4057
rect 4500 -10482 4534 4057
rect 4534 -10482 4539 4057
rect 5080 -5673 7920 -5607
rect 4873 -6488 5044 -5976
rect 5653 -6602 5702 -5863
rect 6076 -6602 6125 -5865
rect 6504 -6602 6553 -5870
rect 9893 -6002 9956 6358
rect 13341 -6002 13404 6358
rect 16789 -6002 16852 6358
rect 20237 -6002 20300 6358
rect 23685 -6002 23748 6358
rect 27133 -6002 27196 6358
rect 28162 -6188 28169 6530
rect 28169 -6188 28203 6530
rect 28203 -6188 28207 6530
rect 4763 -6879 21770 -6783
rect 22082 -6878 27742 -6782
rect 4496 -10527 4539 -10482
rect 26600 -7051 26958 -6941
rect 4809 -9961 4857 -7994
rect 5410 -9992 5454 -9014
rect 8454 -9958 8497 -7988
rect 8577 -9188 9616 -9136
rect 10217 -9961 10260 -7991
rect 10333 -9961 10376 -7989
rect 12813 -9978 12856 -7989
rect 12929 -9963 12972 -7985
rect 15077 -9978 15120 -7987
rect 17151 -9958 17194 -7983
rect 19295 -9955 19338 -7985
rect 21449 -9949 21492 -7985
rect 23593 -9949 23636 -7985
rect 25808 -9966 25851 -7987
rect 4763 -10256 27915 -10161
rect 4595 -10569 28143 -10550
rect 28143 -10569 28200 -10550
rect 4595 -10595 28200 -10569
rect 28361 -10618 28405 6778
rect 28405 -10618 28408 6778
rect 4386 -10741 28323 -10704
rect 4386 -10752 28323 -10741
<< metal1 >>
rect 4253 6871 28439 6899
rect 4253 6817 4427 6871
rect 28261 6817 28439 6871
rect 4253 6786 28439 6817
rect 4253 6767 4356 6786
rect 4253 -10614 4270 6767
rect 4320 6319 4356 6767
rect 28327 6778 28439 6786
rect 9650 6644 28223 6656
rect 9650 6594 9678 6644
rect 28150 6594 28223 6644
rect 9650 6579 28223 6594
rect 28149 6530 28223 6579
rect 9713 6433 27364 6511
rect 4320 6306 4480 6319
rect 4320 6295 8702 6306
rect 4320 6207 6886 6295
rect 7400 6207 8702 6295
rect 4320 6197 8702 6207
rect 4320 6171 4480 6197
rect 4320 4793 4356 6171
rect 6087 5973 6255 5990
rect 6087 5872 6108 5973
rect 6233 5872 6255 5973
rect 6087 5856 6255 5872
rect 8199 5973 8367 5990
rect 8199 5872 8220 5973
rect 8345 5872 8367 5973
rect 8199 5856 8367 5872
rect 6253 5635 6807 5692
rect 8682 5591 9637 5607
rect 8682 5584 9510 5591
rect 4477 5389 9510 5584
rect 8682 5357 9510 5389
rect 4466 5261 4537 5274
rect 4466 4869 4475 5261
rect 4528 4869 4537 5261
rect 4466 4856 4537 4869
rect 6576 5266 6647 5280
rect 6576 4876 6587 5266
rect 6636 4876 6647 5266
rect 9489 5204 9510 5357
rect 9622 5204 9637 5591
rect 9489 5188 9637 5204
rect 6576 4862 6647 4876
rect 4320 4758 4479 4793
rect 4320 4744 8701 4758
rect 4320 4664 6887 4744
rect 4320 4645 4479 4664
rect 7401 4664 8701 4744
rect 4320 -10614 4356 4645
rect 4481 4143 9617 4159
rect 4481 4126 4582 4143
rect 4481 -10527 4496 4126
rect 4539 4098 4582 4126
rect 9580 4098 9617 4143
rect 4539 4075 9617 4098
rect 4539 -6592 4552 4075
rect 8857 3720 9398 3734
rect 8857 3711 8876 3720
rect 5119 3474 5551 3710
rect 7519 3640 8876 3711
rect 8857 3632 8876 3640
rect 9379 3632 9398 3720
rect 8857 3619 9398 3632
rect 5119 3142 5551 3378
rect 7519 3308 7951 3545
rect 5119 2810 5551 3046
rect 7519 2976 7951 3213
rect 5119 2478 5551 2714
rect 7519 2644 7951 2881
rect 5119 2146 5551 2382
rect 7519 2312 7951 2549
rect 5119 1814 5551 2050
rect 7519 1980 7951 2217
rect 5119 1482 5551 1718
rect 7519 1648 7951 1885
rect 5119 1150 5551 1386
rect 7519 1316 7951 1553
rect 5119 818 5551 1054
rect 7519 984 7951 1221
rect 7519 657 7951 889
rect 8426 657 8476 659
rect 7519 607 8476 657
rect 5117 181 5549 417
rect 7519 347 7951 607
rect 5117 -151 5549 85
rect 7517 15 7949 252
rect 5117 -483 5549 -247
rect 7517 -317 7949 -80
rect 5117 -815 5549 -579
rect 7517 -649 7949 -412
rect 5117 -1147 5549 -911
rect 7517 -981 7949 -744
rect 5117 -1479 5549 -1243
rect 7517 -1313 7949 -1076
rect 5117 -1811 5549 -1575
rect 7517 -1645 7949 -1408
rect 5117 -2143 5549 -1907
rect 7517 -1977 7949 -1740
rect 5117 -2475 5549 -2239
rect 7517 -2309 7949 -2072
rect 5117 -2807 5549 -2571
rect 7517 -2641 7949 -2404
rect 5117 -3139 5549 -2903
rect 7517 -2973 7949 -2736
rect 5117 -3471 5549 -3235
rect 7517 -3305 7949 -3068
rect 5117 -3803 5549 -3567
rect 7517 -3637 7949 -3400
rect 5117 -4135 5549 -3899
rect 7517 -3969 7949 -3732
rect 5117 -4467 5549 -4231
rect 7517 -4301 7949 -4064
rect 5117 -4799 5549 -4563
rect 7517 -4633 7949 -4396
rect 5117 -5131 5549 -4895
rect 7517 -4965 7949 -4728
rect 5117 -5463 5549 -5227
rect 7517 -5297 7949 -5060
rect 7517 -5560 7949 -5392
rect 5047 -5561 8199 -5560
rect 4854 -5607 8199 -5561
rect 4854 -5673 5080 -5607
rect 7920 -5673 8199 -5607
rect 4854 -5686 8199 -5673
rect 4854 -5954 5063 -5686
rect 7517 -5688 7949 -5686
rect 5432 -5804 6755 -5772
rect 5628 -5863 5724 -5850
rect 4855 -5976 5062 -5954
rect 4855 -6488 4873 -5976
rect 5044 -6488 5062 -5976
rect 4855 -6504 5062 -6488
rect 5628 -6592 5653 -5863
rect 4539 -6602 5653 -6592
rect 5702 -6108 5724 -5863
rect 6049 -5865 6145 -5850
rect 5702 -6284 5802 -6108
rect 5702 -6592 5724 -6284
rect 5870 -6381 5904 -6024
rect 6049 -6592 6076 -5865
rect 5702 -6602 6076 -6592
rect 6125 -6106 6145 -5865
rect 6479 -5870 6575 -5850
rect 6125 -6282 6230 -6106
rect 6125 -6592 6145 -6282
rect 6297 -6375 6331 -6018
rect 6479 -6592 6504 -5870
rect 6125 -6602 6504 -6592
rect 6553 -6113 6575 -5870
rect 6553 -6289 6656 -6113
rect 6553 -6592 6575 -6289
rect 6721 -6375 6755 -5804
rect 6816 -6457 6871 -6092
rect 8426 -6405 8476 607
rect 9713 -6102 9791 6433
rect 9870 6358 9989 6395
rect 9870 -5864 9893 6358
rect 9956 -5864 9989 6358
rect 9870 -6026 9880 -5864
rect 9980 -6026 9989 -5864
rect 9870 -6035 9989 -6026
rect 10143 -6102 10174 6433
rect 10301 -6102 10332 6433
rect 10459 -6102 10490 6433
rect 10617 -6102 10648 6433
rect 10775 -6102 10806 6433
rect 10933 -6102 10964 6433
rect 11091 -6102 11122 6433
rect 11249 -6102 11280 6433
rect 11407 -6102 11438 6433
rect 11565 -6102 11596 6433
rect 11723 -6102 11754 6433
rect 11881 -6102 11912 6433
rect 12039 -6102 12070 6433
rect 12197 -6102 12228 6433
rect 12355 -6102 12386 6433
rect 12513 -6102 12544 6433
rect 12671 -6102 12702 6433
rect 12829 -6102 12860 6433
rect 12987 -6102 13018 6433
rect 13145 -6102 13176 6433
rect 13318 6358 13437 6395
rect 13318 -5864 13341 6358
rect 13404 -5864 13437 6358
rect 13318 -6026 13328 -5864
rect 13428 -6026 13437 -5864
rect 13318 -6035 13437 -6026
rect 13591 -6102 13622 6433
rect 13749 -6102 13780 6433
rect 13907 -6102 13938 6433
rect 14065 -6102 14096 6433
rect 14223 -6102 14254 6433
rect 14381 -6102 14412 6433
rect 14539 -6102 14570 6433
rect 14697 -6102 14728 6433
rect 14855 -6102 14886 6433
rect 15013 -6102 15044 6433
rect 15171 -6102 15202 6433
rect 15329 -6102 15360 6433
rect 15487 -6102 15518 6433
rect 15645 -6102 15676 6433
rect 15803 -6102 15834 6433
rect 15961 -6102 15992 6433
rect 16119 -6102 16150 6433
rect 16277 -6102 16308 6433
rect 16435 -6102 16466 6433
rect 16593 -6102 16624 6433
rect 16766 6358 16885 6395
rect 16766 -5864 16789 6358
rect 16852 -5864 16885 6358
rect 16766 -6026 16776 -5864
rect 16876 -6026 16885 -5864
rect 16766 -6035 16885 -6026
rect 17039 -6102 17070 6433
rect 17197 -6102 17228 6433
rect 17355 -6102 17386 6433
rect 17513 -6102 17544 6433
rect 17671 -6102 17702 6433
rect 17829 -6102 17860 6433
rect 17987 -6102 18018 6433
rect 18145 -6102 18176 6433
rect 18303 -6102 18334 6433
rect 18461 -6102 18492 6433
rect 18619 -6102 18650 6433
rect 18777 -6102 18808 6433
rect 18935 -6102 18966 6433
rect 19093 -6102 19124 6433
rect 19251 -6102 19282 6433
rect 19409 -6102 19440 6433
rect 19567 -6102 19598 6433
rect 19725 -6102 19756 6433
rect 19883 -6102 19914 6433
rect 20041 -6102 20072 6433
rect 20214 6358 20333 6395
rect 20214 -5864 20237 6358
rect 20300 -5864 20333 6358
rect 20214 -6026 20224 -5864
rect 20324 -6026 20333 -5864
rect 20214 -6035 20333 -6026
rect 20487 -6102 20518 6433
rect 20645 -6102 20676 6433
rect 20803 -6102 20834 6433
rect 20961 -6102 20992 6433
rect 21119 -6102 21150 6433
rect 21277 -6102 21308 6433
rect 21435 -6102 21466 6433
rect 21593 -6102 21624 6433
rect 21751 -6102 21782 6433
rect 21909 -6102 21940 6433
rect 22067 -6102 22098 6433
rect 22225 -6102 22256 6433
rect 22383 -6102 22414 6433
rect 22541 -6102 22572 6433
rect 22699 -6102 22730 6433
rect 22857 -6102 22888 6433
rect 23015 -6102 23046 6433
rect 23173 -6102 23204 6433
rect 23331 -6102 23362 6433
rect 23489 -6102 23520 6433
rect 23662 6358 23781 6395
rect 23662 -5864 23685 6358
rect 23748 -5864 23781 6358
rect 23662 -6026 23672 -5864
rect 23772 -6026 23781 -5864
rect 23662 -6035 23781 -6026
rect 23935 -6102 23966 6433
rect 24093 -6102 24124 6433
rect 24251 -6102 24282 6433
rect 24409 -6102 24440 6433
rect 24567 -6102 24598 6433
rect 24725 -6102 24756 6433
rect 24883 -6102 24914 6433
rect 25041 -6102 25072 6433
rect 25199 -6102 25230 6433
rect 25357 -6102 25388 6433
rect 25515 -6102 25546 6433
rect 25673 -6102 25704 6433
rect 25831 -6102 25862 6433
rect 25989 -6102 26020 6433
rect 26147 -6102 26178 6433
rect 26305 -6102 26336 6433
rect 26463 -6102 26494 6433
rect 26621 -6102 26652 6433
rect 26779 -6102 26810 6433
rect 26937 -6102 26968 6433
rect 27110 6358 27229 6395
rect 27110 -5864 27133 6358
rect 27196 -5864 27229 6358
rect 27110 -6026 27120 -5864
rect 27220 -6026 27229 -5864
rect 27110 -6035 27229 -6026
rect 27286 -6102 27364 6433
rect 9713 -6180 27364 -6102
rect 10699 -6194 10917 -6180
rect 10699 -6386 10717 -6194
rect 10901 -6386 10917 -6194
rect 10699 -6398 10917 -6386
rect 28149 -6188 28162 6530
rect 28207 -6188 28223 6530
rect 10699 -6404 10916 -6398
rect 6816 -6512 27345 -6457
rect 28149 -6536 28223 -6188
rect 6553 -6602 21891 -6592
rect 4539 -6605 21891 -6602
rect 4539 -6606 9393 -6605
rect 4539 -6783 4854 -6606
rect 5250 -6783 9393 -6606
rect 9707 -6783 21891 -6605
rect 4539 -6879 4763 -6783
rect 21770 -6879 21891 -6783
rect 4539 -6909 4854 -6879
rect 5250 -6909 9393 -6879
rect 4539 -6917 9393 -6909
rect 9707 -6917 21891 -6879
rect 4539 -6927 21891 -6917
rect 22029 -6605 28260 -6592
rect 22029 -6782 23670 -6605
rect 23768 -6782 27118 -6605
rect 27216 -6782 28260 -6605
rect 22029 -6878 22082 -6782
rect 27742 -6878 28260 -6782
rect 22029 -6915 23670 -6878
rect 23768 -6915 27118 -6878
rect 27216 -6915 28260 -6878
rect 22029 -6927 28260 -6915
rect 4539 -10527 4552 -6927
rect 4789 -7552 4903 -6927
rect 5599 -7422 5708 -7068
rect 6363 -7344 6646 -7166
rect 6018 -7823 6049 -7687
rect 6263 -7757 6294 -7677
rect 6485 -7689 6524 -7344
rect 6702 -7420 6734 -7078
rect 6805 -7612 6847 -7147
rect 6932 -7556 7060 -6927
rect 7726 -7427 7827 -7076
rect 8525 -7341 8789 -7164
rect 6805 -7654 8536 -7612
rect 6485 -7728 7581 -7689
rect 8639 -7701 8678 -7341
rect 8852 -7415 8884 -7073
rect 8956 -7614 8998 -7152
rect 9081 -7533 9208 -6927
rect 9887 -7422 9988 -7071
rect 10675 -7168 10939 -7157
rect 10675 -7321 10716 -7168
rect 10904 -7321 10939 -7168
rect 10675 -7334 10939 -7321
rect 10998 -7614 11039 -7090
rect 8956 -7655 11039 -7614
rect 6263 -7788 7157 -7757
rect 4776 -7843 4917 -7841
rect 4776 -7994 4919 -7843
rect 6007 -7854 7083 -7823
rect 4776 -9961 4809 -7994
rect 4857 -8841 4919 -7994
rect 5791 -8701 5875 -7974
rect 7052 -8561 7083 -7854
rect 6926 -8592 7083 -8561
rect 6926 -8789 6957 -8592
rect 7126 -8635 7157 -7788
rect 7435 -8482 7469 -7976
rect 7542 -8427 7581 -7728
rect 7875 -8480 7921 -7708
rect 7988 -7740 8678 -7701
rect 7988 -8432 8027 -7740
rect 8864 -7784 10052 -7739
rect 8408 -7988 8557 -7848
rect 9998 -7962 10052 -7784
rect 5714 -8820 6957 -8789
rect 6999 -8666 7157 -8635
rect 4857 -9961 4917 -8841
rect 4776 -10088 4917 -9961
rect 5379 -9014 5535 -8987
rect 5379 -9375 5410 -9014
rect 5454 -9375 5535 -9014
rect 5379 -9577 5397 -9375
rect 5520 -9577 5535 -9375
rect 5379 -9992 5410 -9577
rect 5454 -9992 5535 -9577
rect 5574 -9747 5645 -9261
rect 5379 -10018 5535 -9992
rect 5714 -9977 5745 -8820
rect 6999 -8892 7030 -8666
rect 7426 -8707 7472 -8482
rect 6140 -8923 7030 -8892
rect 7078 -8761 7709 -8707
rect 5811 -9890 5846 -9270
rect 5997 -9754 6068 -9260
rect 6140 -9797 6171 -8923
rect 6556 -9014 6937 -8993
rect 6556 -9168 6595 -9014
rect 6909 -9092 6937 -9014
rect 7078 -9092 7132 -8761
rect 6909 -9146 7132 -9092
rect 6909 -9168 6937 -9146
rect 6556 -9191 6937 -9168
rect 7323 -9258 7369 -8913
rect 7440 -9313 7470 -8998
rect 7640 -9075 7709 -8761
rect 7531 -9256 7822 -9075
rect 7887 -9294 7917 -9012
rect 7976 -9255 8306 -9073
rect 7440 -9414 7470 -9347
rect 6235 -9455 7817 -9414
rect 6419 -9541 7712 -9490
rect 6231 -9747 6235 -9696
rect 6419 -9797 6470 -9541
rect 6111 -9848 6470 -9797
rect 6551 -9699 7398 -9657
rect 6551 -9890 6593 -9699
rect 5811 -9932 6593 -9890
rect 7437 -9891 7474 -9604
rect 6637 -9911 7474 -9891
rect 6637 -9930 7442 -9911
rect 6637 -9977 6676 -9930
rect 5714 -10020 6678 -9977
rect 7544 -10088 7598 -9657
rect 7675 -9890 7712 -9541
rect 7776 -9851 7817 -9455
rect 7881 -9890 7918 -9294
rect 7675 -9906 7918 -9890
rect 7675 -9927 7884 -9906
rect 7985 -10088 8039 -9657
rect 8243 -9707 8306 -9255
rect 8408 -9958 8454 -7988
rect 8497 -9080 8557 -7988
rect 9220 -8899 9312 -7982
rect 9990 -8008 10052 -7962
rect 9998 -8239 10052 -8008
rect 10081 -8559 10124 -7655
rect 11103 -7707 11145 -7149
rect 11223 -7558 11360 -6927
rect 12048 -7416 12140 -7070
rect 12825 -7617 12893 -7146
rect 12952 -7549 13087 -6927
rect 14064 -7430 14156 -7084
rect 10297 -7749 11145 -7707
rect 11556 -7685 12893 -7617
rect 14071 -7587 14141 -7430
rect 15149 -7587 15219 -7137
rect 15286 -7550 15412 -6927
rect 16104 -7420 16196 -7074
rect 16878 -7330 17144 -7160
rect 17208 -7412 17240 -7078
rect 14071 -7657 15219 -7587
rect 10297 -7791 10427 -7749
rect 10028 -8602 10124 -8559
rect 10155 -7989 10427 -7791
rect 11556 -7977 11624 -7685
rect 10155 -7991 10333 -7989
rect 8497 -9136 9665 -9080
rect 10028 -9093 10071 -8602
rect 10155 -9044 10217 -7991
rect 8497 -9188 8577 -9136
rect 9616 -9188 9665 -9136
rect 8497 -9253 9665 -9188
rect 9905 -9136 10071 -9093
rect 8497 -9958 8557 -9253
rect 8678 -9515 8774 -9253
rect 8902 -9457 8930 -9440
rect 8677 -9695 8847 -9515
rect 8408 -10088 8557 -9958
rect 8902 -9962 8930 -9467
rect 9121 -9515 9217 -9253
rect 9345 -9457 9373 -9440
rect 9121 -9696 9302 -9515
rect 9345 -9962 9373 -9467
rect 9566 -9515 9662 -9253
rect 9566 -9679 9746 -9515
rect 9567 -9696 9746 -9679
rect 9792 -9962 9820 -9439
rect 9905 -9709 9948 -9136
rect 10158 -9280 10217 -9044
rect 8902 -9990 9820 -9962
rect 10155 -9961 10217 -9280
rect 10260 -9961 10333 -7991
rect 10376 -9016 10427 -7989
rect 10488 -8825 10558 -8041
rect 10376 -9019 10480 -9016
rect 10376 -9589 10557 -9019
rect 11533 -9475 11644 -7977
rect 12629 -8234 12697 -7685
rect 12764 -7842 12894 -7816
rect 12764 -7985 13018 -7842
rect 12764 -7989 12929 -7985
rect 12626 -9400 12696 -8616
rect 12764 -9589 12813 -7989
rect 10376 -9773 12813 -9589
rect 10376 -9961 10557 -9773
rect 10155 -10088 10557 -9961
rect 12764 -9978 12813 -9773
rect 12856 -9963 12929 -7989
rect 12972 -9963 13018 -7985
rect 12856 -9978 13018 -9963
rect 13844 -9973 13994 -7972
rect 14896 -9896 14966 -7657
rect 17308 -7730 17360 -7148
rect 17440 -7556 17566 -6927
rect 18242 -7422 18334 -7076
rect 19028 -7338 19294 -7168
rect 19364 -7416 19396 -7082
rect 16116 -7786 17360 -7730
rect 18248 -7730 18304 -7422
rect 19464 -7730 19510 -7154
rect 19584 -7548 19716 -6927
rect 26562 -6941 26994 -6927
rect 26562 -7051 26600 -6941
rect 26958 -7051 26994 -6941
rect 19904 -7418 19996 -7072
rect 20184 -7334 20446 -7164
rect 20160 -7388 20206 -7336
rect 20142 -7434 20206 -7388
rect 20638 -7426 20730 -7080
rect 20910 -7332 21172 -7162
rect 20886 -7388 20932 -7338
rect 20868 -7434 20932 -7388
rect 21356 -7426 21448 -7080
rect 21639 -7388 21685 -7153
rect 21592 -7434 21685 -7388
rect 21639 -7601 21685 -7434
rect 22164 -7435 22595 -7200
rect 26562 -7268 26994 -7051
rect 27433 -7535 27477 -7150
rect 27548 -7601 27580 -7084
rect 21639 -7647 27818 -7601
rect 18248 -7786 25676 -7730
rect 15034 -7987 15164 -7848
rect 16116 -7934 16172 -7786
rect 12764 -10088 13018 -9978
rect 15034 -9978 15077 -7987
rect 15120 -9978 15164 -7987
rect 16063 -9977 16213 -7976
rect 17038 -9894 17094 -7786
rect 17131 -7983 17217 -7834
rect 17131 -9958 17151 -7983
rect 17194 -9958 17217 -7983
rect 15034 -10088 15164 -9978
rect 17131 -10088 17217 -9958
rect 17248 -8313 17314 -8030
rect 17248 -8731 17314 -8377
rect 17248 -9149 17314 -8795
rect 17248 -9567 17314 -9213
rect 17248 -9985 17314 -9631
rect 18201 -9973 18351 -7972
rect 19184 -9904 19240 -7786
rect 19277 -7985 19363 -7841
rect 19277 -9955 19295 -7985
rect 19338 -9955 19363 -7985
rect 17248 -10056 17314 -10049
rect 19277 -10088 19363 -9955
rect 19394 -8313 19460 -8030
rect 19394 -8731 19460 -8377
rect 19394 -9149 19460 -8795
rect 19394 -9567 19460 -9213
rect 19394 -9985 19460 -9631
rect 20328 -9966 20478 -7965
rect 21336 -9900 21392 -7786
rect 21426 -7985 21512 -7841
rect 21426 -9949 21449 -7985
rect 21492 -9949 21512 -7985
rect 19394 -10056 19460 -10049
rect 21426 -10088 21512 -9949
rect 21540 -8313 21606 -8030
rect 21540 -8731 21606 -8377
rect 21540 -9149 21606 -8795
rect 21540 -9567 21606 -9213
rect 21540 -9985 21606 -9631
rect 22428 -9966 22578 -7965
rect 23478 -9900 23534 -7786
rect 23572 -7985 23658 -7836
rect 23572 -9949 23593 -7985
rect 23636 -9949 23658 -7985
rect 21540 -10056 21606 -10049
rect 23572 -10088 23658 -9949
rect 23686 -8313 23752 -8030
rect 23686 -8731 23752 -8377
rect 23686 -9149 23752 -8795
rect 23686 -9567 23752 -9213
rect 23686 -9985 23752 -9631
rect 24596 -9970 24746 -7969
rect 25620 -9884 25676 -7786
rect 25772 -7987 25896 -7838
rect 25772 -9966 25808 -7987
rect 25851 -9966 25896 -7987
rect 26758 -9966 26908 -7965
rect 27772 -9908 27818 -7647
rect 27868 -8313 27935 -7370
rect 27934 -8377 27935 -8313
rect 27868 -8731 27935 -8377
rect 27934 -8795 27935 -8731
rect 27868 -9149 27935 -8795
rect 27934 -9213 27935 -9149
rect 27868 -9567 27935 -9213
rect 27934 -9631 27935 -9567
rect 23686 -10056 23752 -10049
rect 25772 -10088 25896 -9966
rect 27868 -9985 27935 -9631
rect 27934 -10049 27935 -9985
rect 27868 -10055 27935 -10049
rect 27993 -10088 28260 -6927
rect 4690 -10161 28260 -10088
rect 4690 -10256 4763 -10161
rect 27915 -10256 28260 -10161
rect 4690 -10474 4991 -10256
rect 5513 -10288 28260 -10256
rect 5513 -10364 5664 -10288
rect 8150 -10290 28260 -10288
rect 8150 -10355 8406 -10290
rect 27898 -10355 28260 -10290
rect 8150 -10364 28260 -10355
rect 5513 -10474 28260 -10364
rect 4690 -10483 28260 -10474
rect 4481 -10530 4552 -10527
rect 4481 -10550 28227 -10530
rect 4481 -10595 4595 -10550
rect 28200 -10595 28227 -10550
rect 4481 -10613 28227 -10595
rect 4253 -10665 4356 -10614
rect 28327 -10618 28361 6778
rect 28408 -10618 28439 6778
rect 28327 -10665 28439 -10618
rect 4253 -10704 28439 -10665
rect 4253 -10752 4386 -10704
rect 28323 -10752 28439 -10704
rect 4253 -10775 28439 -10752
<< via1 >>
rect 6886 6207 7400 6295
rect 4780 5635 5319 5692
rect 9510 5204 9622 5591
rect 6887 4656 7401 4744
rect 8876 3632 9379 3720
rect 4873 -6488 5044 -5976
rect 9880 -6002 9893 -5864
rect 9893 -6002 9956 -5864
rect 9956 -6002 9980 -5864
rect 9880 -6026 9980 -6002
rect 13328 -6002 13341 -5864
rect 13341 -6002 13404 -5864
rect 13404 -6002 13428 -5864
rect 13328 -6026 13428 -6002
rect 16776 -6002 16789 -5864
rect 16789 -6002 16852 -5864
rect 16852 -6002 16876 -5864
rect 16776 -6026 16876 -6002
rect 20224 -6002 20237 -5864
rect 20237 -6002 20300 -5864
rect 20300 -6002 20324 -5864
rect 20224 -6026 20324 -6002
rect 23672 -6002 23685 -5864
rect 23685 -6002 23748 -5864
rect 23748 -6002 23772 -5864
rect 23672 -6026 23772 -6002
rect 27120 -6002 27133 -5864
rect 27133 -6002 27196 -5864
rect 27196 -6002 27220 -5864
rect 27120 -6026 27220 -6002
rect 10717 -6386 10901 -6194
rect 4854 -6783 5250 -6606
rect 9393 -6783 9707 -6605
rect 4854 -6879 5250 -6783
rect 9393 -6879 9707 -6783
rect 4854 -6909 5250 -6879
rect 9393 -6917 9707 -6879
rect 23670 -6782 23768 -6605
rect 27118 -6782 27216 -6605
rect 23670 -6878 23768 -6782
rect 27118 -6878 27216 -6782
rect 23670 -6915 23768 -6878
rect 27118 -6915 27216 -6878
rect 10716 -7321 10904 -7168
rect 5397 -9577 5410 -9375
rect 5410 -9577 5454 -9375
rect 5454 -9577 5520 -9375
rect 6595 -9168 6909 -9014
rect 17248 -8377 17314 -8313
rect 17248 -8795 17314 -8731
rect 17248 -9213 17314 -9149
rect 17248 -9631 17314 -9567
rect 17248 -10049 17314 -9985
rect 19394 -8377 19460 -8313
rect 19394 -8795 19460 -8731
rect 19394 -9213 19460 -9149
rect 19394 -9631 19460 -9567
rect 19394 -10049 19460 -9985
rect 21540 -8377 21606 -8313
rect 21540 -8795 21606 -8731
rect 21540 -9213 21606 -9149
rect 21540 -9631 21606 -9567
rect 21540 -10049 21606 -9985
rect 23686 -8377 23752 -8313
rect 23686 -8795 23752 -8731
rect 23686 -9213 23752 -9149
rect 23686 -9631 23752 -9567
rect 27868 -8377 27934 -8313
rect 27868 -8795 27934 -8731
rect 27868 -9213 27934 -9149
rect 27868 -9631 27934 -9567
rect 23686 -10049 23752 -9985
rect 27868 -10049 27934 -9985
rect 4991 -10256 5513 -10235
rect 4991 -10474 5513 -10256
rect 5664 -10364 8150 -10288
rect 8406 -10355 27898 -10290
<< metal2 >>
rect 4779 5692 5319 6899
rect 6055 6695 6255 6895
rect 7058 6892 7258 6893
rect 6130 5974 6187 6695
rect 6871 6295 7411 6892
rect 8169 6695 8369 6895
rect 6871 6207 6886 6295
rect 7400 6207 7411 6295
rect 4779 5635 4780 5692
rect 4473 4430 4529 4944
rect 4779 4640 5319 5635
rect 6585 4436 6641 4983
rect 6871 4744 7411 6207
rect 8237 5976 8294 6695
rect 8806 6089 9443 6867
rect 27522 6392 28159 6500
rect 6871 4656 6887 4744
rect 7401 4656 7411 4744
rect 6871 4633 7411 4656
rect 8806 5689 27440 6089
rect 8806 4871 9443 5689
rect 9499 5591 9637 5607
rect 9499 5204 9510 5591
rect 9622 5589 9637 5591
rect 27522 5589 27645 6392
rect 9622 5204 27645 5589
rect 9499 5189 27645 5204
rect 9499 5188 9637 5189
rect 8806 4471 27440 4871
rect 4473 4374 6286 4430
rect 6585 4380 6715 4436
rect 4701 -5813 5341 -5767
rect 4701 -9651 4747 -5813
rect 4855 -5976 5062 -5954
rect 4855 -6488 4873 -5976
rect 5044 -6488 5062 -5976
rect 4855 -6504 5062 -6488
rect 5373 -5986 6010 -5944
rect 4842 -6606 5263 -6588
rect 4842 -6909 4854 -6606
rect 5250 -6909 5263 -6606
rect 4842 -6927 5263 -6909
rect 4842 -9360 4996 -6927
rect 5373 -6960 5415 -5986
rect 5968 -6297 6010 -5986
rect 6230 -6357 6286 4374
rect 6185 -6375 6328 -6357
rect 6185 -6422 6205 -6375
rect 5871 -6471 6205 -6422
rect 6185 -6623 6205 -6471
rect 6303 -6623 6328 -6375
rect 6185 -6644 6328 -6623
rect 5046 -7002 5415 -6960
rect 5046 -7392 5088 -7002
rect 6395 -7040 6439 -6274
rect 6659 -6557 6715 4380
rect 8806 3720 9443 4471
rect 27522 4371 27645 5189
rect 9867 3971 27645 4371
rect 8806 3632 8876 3720
rect 9379 3653 9443 3720
rect 9379 3632 27440 3653
rect 8806 3253 27440 3632
rect 8806 2435 9443 3253
rect 27522 3153 27645 3971
rect 9867 2753 27645 3153
rect 8806 2035 27440 2435
rect 8806 1217 9443 2035
rect 27522 1935 27645 2753
rect 9867 1535 27645 1935
rect 8806 817 27440 1217
rect 8806 -1 9443 817
rect 27522 717 27645 1535
rect 9867 317 27645 717
rect 8806 -401 27440 -1
rect 8806 -1219 9443 -401
rect 27522 -501 27645 317
rect 9867 -901 27645 -501
rect 8806 -1619 27440 -1219
rect 8806 -2437 9443 -1619
rect 27522 -1719 27645 -901
rect 9867 -2119 27645 -1719
rect 8806 -2837 27440 -2437
rect 8806 -3655 9443 -2837
rect 27522 -2937 27645 -2119
rect 9867 -3337 27645 -2937
rect 8806 -4055 27440 -3655
rect 8806 -4873 9443 -4055
rect 27522 -4155 27645 -3337
rect 9867 -4555 27645 -4155
rect 8806 -5273 27440 -4873
rect 8806 -5990 9443 -5273
rect 27522 -5373 27645 -4555
rect 9867 -5773 27645 -5373
rect 9869 -5864 9989 -5852
rect 9869 -6026 9880 -5864
rect 9980 -6026 9989 -5864
rect 8418 -6554 8480 -6402
rect 6619 -6574 6762 -6557
rect 6619 -6822 6643 -6574
rect 6741 -6822 6762 -6574
rect 8296 -6567 8593 -6554
rect 8296 -6642 8311 -6567
rect 8577 -6642 8593 -6567
rect 8296 -6654 8593 -6642
rect 9378 -6605 9726 -6588
rect 6619 -6844 6762 -6822
rect 9378 -6917 9393 -6605
rect 9707 -6917 9726 -6605
rect 9378 -6931 9726 -6917
rect 9869 -6592 9989 -6026
rect 13317 -5864 13437 -5852
rect 13317 -6026 13328 -5864
rect 13428 -6026 13437 -5864
rect 10699 -6194 10916 -6184
rect 10699 -6386 10717 -6194
rect 10901 -6386 10916 -6194
rect 10699 -6404 10916 -6386
rect 13317 -6592 13437 -6026
rect 16765 -5864 16885 -5852
rect 16765 -6026 16776 -5864
rect 16876 -6026 16885 -5864
rect 16765 -6592 16885 -6026
rect 20213 -5864 20333 -5852
rect 20213 -6026 20224 -5864
rect 20324 -6026 20333 -5864
rect 20213 -6592 20333 -6026
rect 23661 -5864 23781 -5852
rect 23661 -6026 23672 -5864
rect 23772 -6026 23781 -5864
rect 23661 -6592 23781 -6026
rect 27109 -5864 27229 -5852
rect 27109 -6026 27120 -5864
rect 27220 -6026 27229 -5864
rect 27522 -5877 27645 -5773
rect 28052 -5877 28159 6392
rect 27522 -6009 28159 -5877
rect 27109 -6592 27229 -6026
rect 27307 -6456 27453 -6455
rect 27307 -6512 27703 -6456
rect 27307 -6515 27453 -6512
rect 9869 -6605 27229 -6592
rect 9869 -6915 23670 -6605
rect 23768 -6915 27118 -6605
rect 27216 -6915 27229 -6605
rect 9869 -6925 27229 -6915
rect 5454 -7104 21898 -7040
rect 27647 -7076 27703 -6512
rect 10700 -7168 10913 -7157
rect 10700 -7321 10716 -7168
rect 10904 -7321 10913 -7168
rect 10700 -7334 10913 -7321
rect 5046 -7456 21898 -7392
rect 26640 -7437 27935 -7368
rect 7661 -7511 7912 -7491
rect 5916 -7558 6051 -7539
rect 5916 -7813 5940 -7558
rect 6027 -7813 6051 -7558
rect 6155 -7661 6450 -7642
rect 6155 -7751 6172 -7661
rect 6428 -7751 6450 -7661
rect 7661 -7685 7687 -7511
rect 7891 -7685 7912 -7511
rect 8957 -7517 9235 -7499
rect 8539 -7649 8864 -7610
rect 7661 -7711 7912 -7685
rect 6155 -7777 6450 -7751
rect 8825 -7784 8864 -7649
rect 8957 -7665 8979 -7517
rect 9212 -7665 9235 -7517
rect 8957 -7684 9235 -7665
rect 5916 -7834 6051 -7813
rect 27300 -7895 27363 -7545
rect 5104 -7959 27785 -7895
rect 6784 -8214 8106 -8069
rect 6556 -9014 6937 -8993
rect 6556 -9168 6595 -9014
rect 6909 -9168 6937 -9014
rect 9242 -9071 9281 -7959
rect 12832 -8377 17248 -8313
rect 17314 -8377 19394 -8313
rect 19460 -8377 21540 -8313
rect 21606 -8377 23686 -8313
rect 23752 -8377 27868 -8313
rect 27934 -8377 27944 -8313
rect 12832 -8795 17248 -8731
rect 17314 -8795 19394 -8731
rect 19460 -8795 21540 -8731
rect 21606 -8795 23686 -8731
rect 23752 -8795 27868 -8731
rect 27934 -8795 27944 -8731
rect 6556 -9191 6937 -9168
rect 9008 -9110 9281 -9071
rect 10259 -9087 10344 -9076
rect 7312 -9309 7356 -9203
rect 7312 -9353 8615 -9309
rect 4842 -9375 6334 -9360
rect 4842 -9557 5397 -9375
rect 4843 -9577 5397 -9557
rect 5520 -9577 6334 -9375
rect 4843 -9597 6334 -9577
rect 7024 -9447 8493 -9399
rect 7024 -9651 7070 -9447
rect 4701 -9697 7070 -9651
rect 4965 -10211 5547 -10210
rect 4965 -10235 5548 -10211
rect 4965 -10474 4991 -10235
rect 5513 -10474 5548 -10235
rect 5632 -10288 8179 -10264
rect 5632 -10364 5664 -10288
rect 8150 -10364 8179 -10288
rect 5632 -10382 8179 -10364
rect 4965 -10495 5548 -10474
rect 8240 -10550 8301 -9801
rect 8445 -9945 8493 -9447
rect 8571 -9779 8615 -9353
rect 9008 -9484 9047 -9110
rect 10259 -9215 10270 -9087
rect 9451 -9258 10270 -9215
rect 9451 -9486 9494 -9258
rect 10259 -9304 10270 -9258
rect 10333 -9304 10344 -9087
rect 12832 -9213 17248 -9149
rect 17314 -9213 19394 -9149
rect 19460 -9213 21540 -9149
rect 21606 -9213 23686 -9149
rect 23752 -9213 27868 -9149
rect 27934 -9213 27944 -9149
rect 10259 -9317 10344 -9304
rect 11566 -9779 11610 -9452
rect 12832 -9631 17248 -9567
rect 17314 -9631 19394 -9567
rect 19460 -9631 21540 -9567
rect 21606 -9631 23686 -9567
rect 23752 -9631 27868 -9567
rect 27934 -9631 27944 -9567
rect 8571 -9823 11610 -9779
rect 8445 -9993 9123 -9945
rect 12832 -10049 17248 -9985
rect 17314 -10049 19394 -9985
rect 19460 -10049 21540 -9985
rect 21606 -10049 23686 -9985
rect 23752 -10049 27868 -9985
rect 27934 -10049 27944 -9985
rect 8385 -10290 27916 -10267
rect 8385 -10355 8406 -10290
rect 27898 -10355 27916 -10290
rect 8385 -10370 27916 -10355
rect 8176 -10750 8376 -10550
<< via2 >>
rect 4873 -6488 5044 -5976
rect 6205 -6623 6303 -6375
rect 6643 -6822 6741 -6574
rect 8311 -6642 8577 -6567
rect 9393 -6917 9707 -6605
rect 10717 -6386 10901 -6194
rect 27645 -5877 28052 6392
rect 10716 -7321 10904 -7168
rect 5940 -7813 6027 -7558
rect 6172 -7751 6428 -7661
rect 7687 -7685 7891 -7511
rect 8979 -7665 9212 -7517
rect 6595 -9168 6909 -9014
rect 4991 -10474 5513 -10235
rect 5664 -10364 8150 -10288
rect 10270 -9304 10333 -9087
rect 8406 -10355 27898 -10290
<< metal3 >>
rect 27522 6392 28159 6500
rect 27522 -5877 27645 6392
rect 28052 -5877 28159 6392
rect 4855 -5976 5062 -5954
rect 4855 -6488 4873 -5976
rect 5044 -6488 5062 -5976
rect 8643 -6210 9127 -6191
rect 10699 -6194 10916 -6184
rect 8643 -6306 8665 -6210
rect 9107 -6306 9127 -6210
rect 8643 -6327 9127 -6306
rect 9376 -6230 9726 -6210
rect 4855 -6504 5062 -6488
rect 6185 -6375 6328 -6357
rect 6185 -6623 6205 -6375
rect 6303 -6565 6328 -6375
rect 6303 -6623 6470 -6565
rect 6185 -6644 6470 -6623
rect 6401 -7479 6470 -6644
rect 6619 -6574 6762 -6557
rect 6619 -6806 6643 -6574
rect 5916 -7548 6470 -7479
rect 6547 -6822 6643 -6806
rect 6741 -6822 6762 -6574
rect 6547 -6844 6762 -6822
rect 7764 -6567 8594 -6554
rect 7764 -6619 8311 -6567
rect 6547 -6874 6716 -6844
rect 5916 -7558 6051 -7548
rect 5916 -7813 5940 -7558
rect 6027 -7813 6051 -7558
rect 6547 -7642 6615 -6874
rect 7764 -7491 7830 -6619
rect 8296 -6642 8311 -6619
rect 8577 -6619 8594 -6567
rect 8577 -6642 8593 -6619
rect 8296 -6654 8593 -6642
rect 6155 -7661 6615 -7642
rect 6155 -7751 6172 -7661
rect 6428 -7710 6615 -7661
rect 7661 -7511 7912 -7491
rect 9046 -7499 9126 -6327
rect 9376 -6531 9400 -6230
rect 9705 -6531 9726 -6230
rect 10699 -6386 10717 -6194
rect 10901 -6386 10916 -6194
rect 10699 -6404 10916 -6386
rect 27522 -6228 28159 -5877
rect 9376 -6605 9726 -6531
rect 9376 -6917 9393 -6605
rect 9707 -6917 9726 -6605
rect 9376 -6930 9726 -6917
rect 10700 -7168 10913 -6404
rect 27522 -6539 27540 -6228
rect 28141 -6539 28159 -6228
rect 27522 -6555 28159 -6539
rect 10700 -7321 10716 -7168
rect 10904 -7321 10913 -7168
rect 10700 -7334 10913 -7321
rect 7661 -7685 7687 -7511
rect 7891 -7685 7912 -7511
rect 8957 -7517 9235 -7499
rect 10777 -7504 10841 -7334
rect 8957 -7665 8979 -7517
rect 9212 -7665 9235 -7517
rect 8957 -7684 9235 -7665
rect 10269 -7568 10841 -7504
rect 6428 -7751 6450 -7710
rect 7661 -7711 7912 -7685
rect 6155 -7777 6450 -7751
rect 6328 -7783 6396 -7777
rect 5916 -7834 6051 -7813
rect 6576 -9014 6937 -8993
rect 6576 -9168 6595 -9014
rect 6909 -9168 6937 -9014
rect 10269 -9076 10333 -7568
rect 6576 -9191 6937 -9168
rect 10259 -9087 10344 -9076
rect 10259 -9304 10270 -9087
rect 10333 -9304 10344 -9087
rect 10259 -9317 10344 -9304
rect 4965 -10211 5547 -10210
rect 4965 -10235 5548 -10211
rect 4965 -10474 4991 -10235
rect 5513 -10474 5548 -10235
rect 5632 -10288 8179 -10264
rect 5632 -10364 5664 -10288
rect 8150 -10364 8179 -10288
rect 5632 -10382 8179 -10364
rect 8385 -10290 27916 -10267
rect 8385 -10355 8406 -10290
rect 27898 -10355 27916 -10290
rect 8385 -10370 27916 -10355
rect 4965 -10495 5548 -10474
<< via3 >>
rect 4873 -6488 5044 -5976
rect 8665 -6306 9107 -6210
rect 9400 -6531 9705 -6230
rect 27540 -6539 28141 -6228
rect 6595 -9168 6909 -9014
rect 4991 -10474 5513 -10235
rect 5664 -10364 8150 -10288
rect 8406 -10355 27898 -10290
<< metal4 >>
rect 4855 -5976 5062 4221
rect 4855 -6488 4873 -5976
rect 5044 -6488 5062 -5976
rect 7812 -5520 8164 2944
rect 7812 -6191 8196 -5520
rect 7812 -6210 9127 -6191
rect 7812 -6306 8665 -6210
rect 9107 -6306 9127 -6210
rect 7812 -6327 9127 -6306
rect 9381 -6228 28395 -6213
rect 9381 -6230 27540 -6228
rect 4855 -10088 5062 -6488
rect 9381 -6531 9400 -6230
rect 9705 -6531 27540 -6230
rect 9381 -6539 27540 -6531
rect 28141 -6539 28395 -6228
rect 9381 -6554 28395 -6539
rect 6556 -9014 6937 -8993
rect 6556 -9069 6595 -9014
rect 6164 -9168 6595 -9069
rect 6909 -9168 6937 -9014
rect 6164 -9189 6937 -9168
rect 6556 -9191 6937 -9189
rect 4291 -10235 28434 -10088
rect 4291 -10474 4991 -10235
rect 5513 -10288 28434 -10235
rect 5513 -10364 5664 -10288
rect 8150 -10290 28434 -10288
rect 8150 -10355 8406 -10290
rect 27898 -10355 28434 -10290
rect 8150 -10364 28434 -10355
rect 5513 -10474 28434 -10364
rect 4291 -10485 28434 -10474
rect 4855 -10495 5548 -10485
use ldo_via_2x2cut  ldo_via_2x2cut_0
timestamp 1717294357
transform 1 0 -10036 0 1 -1046
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_1
timestamp 1717294357
transform 1 0 2638 0 1 -1036
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_2
timestamp 1717294357
transform 1 0 478 0 1 -1034
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_4
timestamp 1717294357
transform 1 0 -7897 0 1 -1044
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_5
timestamp 1717294357
transform 1 0 -10436 0 1 -8
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_6
timestamp 1717294357
transform 1 0 -10855 0 1 -8
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_7
timestamp 1717294357
transform 1 0 -10524 0 1 12348
box 16626 -6492 16764 -6354
use ldo_via_2x2cut  ldo_via_2x2cut_8
timestamp 1717294357
transform 1 0 -8417 0 1 12348
box 16626 -6492 16764 -6354
use ldo_via_4cut  ldo_via_4cut_0
timestamp 1717294357
transform 1 0 4318 0 1 -38
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_1
timestamp 1717294357
transform 1 0 -2166 0 1 -32
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_2
timestamp 1717294357
transform 1 0 46 0 1 -36
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_3
timestamp 1717294357
transform 1 0 -10249 0 1 -48
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_4
timestamp 1717294357
transform -1 0 43520 0 -1 -14383
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_5
timestamp 1717294357
transform 1 0 6418 0 1 -32
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_6
timestamp 1717294357
transform 1 0 8576 0 1 -32
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_7
timestamp 1717294357
transform 1 0 2178 0 1 -36
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_8
timestamp 1717294357
transform 1 0 2206 0 1 832
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_9
timestamp 1717294357
transform 1 0 74 0 1 836
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_10
timestamp 1717294357
transform 1 0 -1974 0 1 474
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_11
timestamp 1717294357
transform 1 0 11258 0 1 366
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_12
timestamp 1717294357
transform 1 0 10693 0 1 495
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_13
timestamp 1717294357
transform 1 0 10746 0 1 -36
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_14
timestamp 1717294357
transform 0 1 35802 -1 0 8578
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_15
timestamp 1717294357
transform 1 0 -4006 0 1 828
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_16
timestamp 1717294357
transform 1 0 -6146 0 1 835
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_17
timestamp 1717294357
transform 0 1 15707 -1 0 7879
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_18
timestamp 1717294357
transform 1 0 -8309 0 1 830
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_19
timestamp 1717294357
transform 0 1 14711 -1 0 7878
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_20
timestamp 1717294357
transform 0 1 15262 -1 0 7879
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_21
timestamp 1717294357
transform 1 0 -10443 0 1 832
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_22
timestamp 1717294357
transform 1 0 -8300 0 1 169
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_23
timestamp 1717294357
transform 1 0 -6990 0 1 269
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_24
timestamp 1717294357
transform 0 1 35574 -1 0 8884
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_25
timestamp 1717294357
transform 0 1 16349 -1 0 9811
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_26
timestamp 1717294357
transform -1 0 25118 0 -1 -17865
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_27
timestamp 1717294357
transform 1 0 -7130 0 1 146
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_28
timestamp 1717294357
transform 0 1 16928 -1 0 6480
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_29
timestamp 1717294357
transform 0 1 17374 -1 0 6476
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_30
timestamp 1717294357
transform 1 0 -7636 0 1 277
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_31
timestamp 1717294357
transform 0 1 13934 -1 0 6605
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_32
timestamp 1717294357
transform 1 0 -9256 0 1 -1774
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_33
timestamp 1717294357
transform 0 1 13513 -1 0 6606
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_34
timestamp 1717294357
transform 0 1 16171 -1 0 6412
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_35
timestamp 1717294357
transform 0 1 15231 -1 0 6957
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_36
timestamp 1717294357
transform -1 0 27686 0 -1 -17384
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_38
timestamp 1717294357
transform -1 0 22382 0 -1 -15654
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_40
timestamp 1717294357
transform 0 1 13928 -1 0 8386
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_41
timestamp 1717294357
transform 1 0 -10768 0 1 2108
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_42
timestamp 1717294357
transform 0 1 14314 -1 0 9906
box 15948 -7932 16222 -7868
use ldo_via_4cut  ldo_via_4cut_43
timestamp 1717294357
transform 0 1 13891 -1 0 9906
box 15948 -7932 16222 -7868
use ldo_via_6cut  ldo_via_6cut_0
timestamp 1717294357
transform 1 0 4049 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1
timestamp 1717294357
transform 1 0 2310 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_2
timestamp 1717294357
transform 1 0 1205 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_3
timestamp 1717294357
transform 1 0 1521 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_4
timestamp 1717294357
transform 1 0 1837 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_5
timestamp 1717294357
transform 1 0 2153 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_6
timestamp 1717294357
transform 1 0 2469 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_7
timestamp 1717294357
transform 1 0 2785 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_8
timestamp 1717294357
transform 1 0 3101 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_9
timestamp 1717294357
transform 1 0 3417 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_10
timestamp 1717294357
transform 1 0 3733 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_11
timestamp 1717294357
transform 1 0 889 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_12
timestamp 1717294357
transform 1 0 1046 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_13
timestamp 1717294357
transform 1 0 1362 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_14
timestamp 1717294357
transform 1 0 1678 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_15
timestamp 1717294357
transform 1 0 1994 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_16
timestamp 1717294357
transform 1 0 2942 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_17
timestamp 1717294357
transform 1 0 2626 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_18
timestamp 1717294357
transform 1 0 3890 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_19
timestamp 1717294357
transform 1 0 3258 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_20
timestamp 1717294357
transform 1 0 3574 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_21
timestamp 1717294357
transform 1 0 3890 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_22
timestamp 1717294357
transform 1 0 3574 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_23
timestamp 1717294357
transform 1 0 3258 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_24
timestamp 1717294357
transform 1 0 2942 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_25
timestamp 1717294357
transform 1 0 2626 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_26
timestamp 1717294357
transform 1 0 2310 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_27
timestamp 1717294357
transform 1 0 1994 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_28
timestamp 1717294357
transform 1 0 1678 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_29
timestamp 1717294357
transform 1 0 1362 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_30
timestamp 1717294357
transform 1 0 1046 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_31
timestamp 1717294357
transform 1 0 4049 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_32
timestamp 1717294357
transform 1 0 3733 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_33
timestamp 1717294357
transform 1 0 3417 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_34
timestamp 1717294357
transform 1 0 3101 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_35
timestamp 1717294357
transform 1 0 2785 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_36
timestamp 1717294357
transform 1 0 2469 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_37
timestamp 1717294357
transform 1 0 2153 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_38
timestamp 1717294357
transform 1 0 1837 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_39
timestamp 1717294357
transform 1 0 1521 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_40
timestamp 1717294357
transform 1 0 1205 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_41
timestamp 1717294357
transform 1 0 889 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_42
timestamp 1717294357
transform 1 0 889 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_43
timestamp 1717294357
transform 1 0 1205 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_44
timestamp 1717294357
transform 1 0 1521 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_45
timestamp 1717294357
transform 1 0 1837 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_46
timestamp 1717294357
transform 1 0 1046 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_47
timestamp 1717294357
transform 1 0 1362 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_48
timestamp 1717294357
transform 1 0 1678 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_49
timestamp 1717294357
transform 1 0 2469 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_50
timestamp 1717294357
transform 1 0 2785 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_51
timestamp 1717294357
transform 1 0 2153 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_52
timestamp 1717294357
transform 1 0 4049 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_53
timestamp 1717294357
transform 1 0 3733 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_54
timestamp 1717294357
transform 1 0 3417 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_55
timestamp 1717294357
transform 1 0 3101 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_56
timestamp 1717294357
transform 1 0 2310 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_57
timestamp 1717294357
transform 1 0 2942 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_58
timestamp 1717294357
transform 1 0 2626 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_59
timestamp 1717294357
transform 1 0 1994 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_60
timestamp 1717294357
transform 1 0 3890 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_61
timestamp 1717294357
transform 1 0 3574 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_62
timestamp 1717294357
transform 1 0 3258 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_63
timestamp 1717294357
transform 1 0 889 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_64
timestamp 1717294357
transform 1 0 1837 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_65
timestamp 1717294357
transform 1 0 1205 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_66
timestamp 1717294357
transform 1 0 1521 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_67
timestamp 1717294357
transform 1 0 1046 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_68
timestamp 1717294357
transform 1 0 1678 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_69
timestamp 1717294357
transform 1 0 1362 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_70
timestamp 1717294357
transform 1 0 2469 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_71
timestamp 1717294357
transform 1 0 2785 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_72
timestamp 1717294357
transform 1 0 2153 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_73
timestamp 1717294357
transform 1 0 4049 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_74
timestamp 1717294357
transform 1 0 3733 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_75
timestamp 1717294357
transform 1 0 3417 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_76
timestamp 1717294357
transform 1 0 3101 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_77
timestamp 1717294357
transform 1 0 2310 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_78
timestamp 1717294357
transform 1 0 2942 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_79
timestamp 1717294357
transform 1 0 2626 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_80
timestamp 1717294357
transform 1 0 1994 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_81
timestamp 1717294357
transform 1 0 3890 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_82
timestamp 1717294357
transform 1 0 3574 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_83
timestamp 1717294357
transform 1 0 3258 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_84
timestamp 1717294357
transform 1 0 889 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_85
timestamp 1717294357
transform 1 0 1837 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_86
timestamp 1717294357
transform 1 0 1205 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_87
timestamp 1717294357
transform 1 0 1521 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_88
timestamp 1717294357
transform 1 0 1046 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_89
timestamp 1717294357
transform 1 0 1678 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_90
timestamp 1717294357
transform 1 0 1362 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_91
timestamp 1717294357
transform 1 0 2469 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_92
timestamp 1717294357
transform 1 0 2785 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_93
timestamp 1717294357
transform 1 0 2153 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_94
timestamp 1717294357
transform 1 0 4049 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_95
timestamp 1717294357
transform 1 0 3733 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_96
timestamp 1717294357
transform 1 0 3417 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_97
timestamp 1717294357
transform 1 0 3101 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_98
timestamp 1717294357
transform 1 0 2310 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_99
timestamp 1717294357
transform 1 0 2942 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_100
timestamp 1717294357
transform 1 0 2626 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_101
timestamp 1717294357
transform 1 0 1994 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_102
timestamp 1717294357
transform 1 0 3890 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_103
timestamp 1717294357
transform 1 0 3574 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_104
timestamp 1717294357
transform 1 0 3258 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_105
timestamp 1717294357
transform 1 0 889 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_106
timestamp 1717294357
transform 1 0 1837 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_107
timestamp 1717294357
transform 1 0 1205 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_108
timestamp 1717294357
transform 1 0 1521 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_109
timestamp 1717294357
transform 1 0 1046 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_110
timestamp 1717294357
transform 1 0 1678 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_111
timestamp 1717294357
transform 1 0 1362 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_112
timestamp 1717294357
transform 1 0 2469 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_113
timestamp 1717294357
transform 1 0 2785 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_114
timestamp 1717294357
transform 1 0 2153 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_115
timestamp 1717294357
transform 1 0 4049 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_116
timestamp 1717294357
transform 1 0 3733 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_117
timestamp 1717294357
transform 1 0 3417 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_118
timestamp 1717294357
transform 1 0 3101 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_119
timestamp 1717294357
transform 1 0 2310 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_120
timestamp 1717294357
transform 1 0 2942 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_121
timestamp 1717294357
transform 1 0 2626 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_122
timestamp 1717294357
transform 1 0 1994 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_123
timestamp 1717294357
transform 1 0 3890 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_124
timestamp 1717294357
transform 1 0 3574 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_125
timestamp 1717294357
transform 1 0 3258 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_126
timestamp 1717294357
transform 1 0 3890 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_127
timestamp 1717294357
transform 1 0 3574 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_128
timestamp 1717294357
transform 1 0 3258 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_129
timestamp 1717294357
transform 1 0 2310 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_130
timestamp 1717294357
transform 1 0 2942 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_131
timestamp 1717294357
transform 1 0 2626 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_132
timestamp 1717294357
transform 1 0 1678 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_133
timestamp 1717294357
transform 1 0 1994 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_134
timestamp 1717294357
transform 1 0 1046 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_135
timestamp 1717294357
transform 1 0 1362 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_136
timestamp 1717294357
transform 1 0 4049 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_137
timestamp 1717294357
transform 1 0 3733 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_138
timestamp 1717294357
transform 1 0 3417 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_139
timestamp 1717294357
transform 1 0 3101 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_140
timestamp 1717294357
transform 1 0 2469 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_141
timestamp 1717294357
transform 1 0 2785 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_142
timestamp 1717294357
transform 1 0 1837 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_143
timestamp 1717294357
transform 1 0 2153 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_144
timestamp 1717294357
transform 1 0 1205 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_145
timestamp 1717294357
transform 1 0 889 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_146
timestamp 1717294357
transform 1 0 1521 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_147
timestamp 1717294357
transform 1 0 1205 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_148
timestamp 1717294357
transform 1 0 889 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_149
timestamp 1717294357
transform 1 0 1837 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_150
timestamp 1717294357
transform 1 0 2153 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_151
timestamp 1717294357
transform 1 0 1521 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_152
timestamp 1717294357
transform 1 0 3417 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_153
timestamp 1717294357
transform 1 0 3101 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_154
timestamp 1717294357
transform 1 0 2469 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_155
timestamp 1717294357
transform 1 0 2785 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_156
timestamp 1717294357
transform 1 0 1046 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_157
timestamp 1717294357
transform 1 0 2310 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_158
timestamp 1717294357
transform 1 0 1678 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_159
timestamp 1717294357
transform 1 0 1994 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_160
timestamp 1717294357
transform 1 0 1362 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_161
timestamp 1717294357
transform 1 0 3258 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_162
timestamp 1717294357
transform 1 0 2942 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_163
timestamp 1717294357
transform 1 0 2626 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_164
timestamp 1717294357
transform 1 0 3733 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_165
timestamp 1717294357
transform 1 0 4049 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_166
timestamp 1717294357
transform 1 0 3574 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_167
timestamp 1717294357
transform 1 0 3890 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_168
timestamp 1717294357
transform 1 0 1205 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_169
timestamp 1717294357
transform 1 0 889 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_170
timestamp 1717294357
transform 1 0 1837 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_171
timestamp 1717294357
transform 1 0 2153 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_172
timestamp 1717294357
transform 1 0 1521 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_173
timestamp 1717294357
transform 1 0 3417 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_174
timestamp 1717294357
transform 1 0 3101 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_175
timestamp 1717294357
transform 1 0 2469 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_176
timestamp 1717294357
transform 1 0 2785 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_177
timestamp 1717294357
transform 1 0 1046 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_178
timestamp 1717294357
transform 1 0 2310 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_179
timestamp 1717294357
transform 1 0 1678 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_180
timestamp 1717294357
transform 1 0 1994 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_181
timestamp 1717294357
transform 1 0 1362 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_182
timestamp 1717294357
transform 1 0 3258 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_183
timestamp 1717294357
transform 1 0 2942 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_184
timestamp 1717294357
transform 1 0 2626 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_185
timestamp 1717294357
transform 1 0 3890 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_186
timestamp 1717294357
transform 1 0 3574 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_187
timestamp 1717294357
transform 1 0 4049 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_188
timestamp 1717294357
transform 1 0 3733 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_189
timestamp 1717294357
transform 1 0 1205 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_190
timestamp 1717294357
transform 1 0 889 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_191
timestamp 1717294357
transform 1 0 1837 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_192
timestamp 1717294357
transform 1 0 2153 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_193
timestamp 1717294357
transform 1 0 1521 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_194
timestamp 1717294357
transform 1 0 3417 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_195
timestamp 1717294357
transform 1 0 3101 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_196
timestamp 1717294357
transform 1 0 2469 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_197
timestamp 1717294357
transform 1 0 2785 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_198
timestamp 1717294357
transform 1 0 4049 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_199
timestamp 1717294357
transform 1 0 3733 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_200
timestamp 1717294357
transform 1 0 3258 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_201
timestamp 1717294357
transform 1 0 2310 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_202
timestamp 1717294357
transform 1 0 2942 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_203
timestamp 1717294357
transform 1 0 2626 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_204
timestamp 1717294357
transform 1 0 1678 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_205
timestamp 1717294357
transform 1 0 1994 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_206
timestamp 1717294357
transform 1 0 1046 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_207
timestamp 1717294357
transform 1 0 1362 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_208
timestamp 1717294357
transform 1 0 7338 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_209
timestamp 1717294357
transform 1 0 7022 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_210
timestamp 1717294357
transform 1 0 5442 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_211
timestamp 1717294357
transform 1 0 5758 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_212
timestamp 1717294357
transform 1 0 6074 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_213
timestamp 1717294357
transform 1 0 4494 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_214
timestamp 1717294357
transform 1 0 5126 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_215
timestamp 1717294357
transform 1 0 4810 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_216
timestamp 1717294357
transform 1 0 6233 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_217
timestamp 1717294357
transform 1 0 5917 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_218
timestamp 1717294357
transform 1 0 5601 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_219
timestamp 1717294357
transform 1 0 4653 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_220
timestamp 1717294357
transform 1 0 5285 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_221
timestamp 1717294357
transform 1 0 4969 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_222
timestamp 1717294357
transform 1 0 4337 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_223
timestamp 1717294357
transform 1 0 7022 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_224
timestamp 1717294357
transform 1 0 7338 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_225
timestamp 1717294357
transform 1 0 6390 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_226
timestamp 1717294357
transform 1 0 6706 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_227
timestamp 1717294357
transform 1 0 7181 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_228
timestamp 1717294357
transform 1 0 7497 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_229
timestamp 1717294357
transform 1 0 6865 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_230
timestamp 1717294357
transform 1 0 6549 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_231
timestamp 1717294357
transform 1 0 4653 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_232
timestamp 1717294357
transform 1 0 4969 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_233
timestamp 1717294357
transform 1 0 4494 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_234
timestamp 1717294357
transform 1 0 4810 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_235
timestamp 1717294357
transform 1 0 4337 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_236
timestamp 1717294357
transform 1 0 4653 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_237
timestamp 1717294357
transform 1 0 4969 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_238
timestamp 1717294357
transform 1 0 4337 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_239
timestamp 1717294357
transform 1 0 4969 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_240
timestamp 1717294357
transform 1 0 4653 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_241
timestamp 1717294357
transform 1 0 4337 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_242
timestamp 1717294357
transform 1 0 4810 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_243
timestamp 1717294357
transform 1 0 4494 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_244
timestamp 1717294357
transform 1 0 4969 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_245
timestamp 1717294357
transform 1 0 4653 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_246
timestamp 1717294357
transform 1 0 4337 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_247
timestamp 1717294357
transform 1 0 4810 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_248
timestamp 1717294357
transform 1 0 4494 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_249
timestamp 1717294357
transform 1 0 4653 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_250
timestamp 1717294357
transform 1 0 4969 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_251
timestamp 1717294357
transform 1 0 4337 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_252
timestamp 1717294357
transform 1 0 4810 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_253
timestamp 1717294357
transform 1 0 4494 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_254
timestamp 1717294357
transform 1 0 4494 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_255
timestamp 1717294357
transform 1 0 4810 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_256
timestamp 1717294357
transform 1 0 7497 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_257
timestamp 1717294357
transform 1 0 7181 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_258
timestamp 1717294357
transform 1 0 7022 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_259
timestamp 1717294357
transform 1 0 7338 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_260
timestamp 1717294357
transform 1 0 6233 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_261
timestamp 1717294357
transform 1 0 6390 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_262
timestamp 1717294357
transform 1 0 6865 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_263
timestamp 1717294357
transform 1 0 6549 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_264
timestamp 1717294357
transform 1 0 6706 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_265
timestamp 1717294357
transform 1 0 5601 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_266
timestamp 1717294357
transform 1 0 5917 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_267
timestamp 1717294357
transform 1 0 5442 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_268
timestamp 1717294357
transform 1 0 5758 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_269
timestamp 1717294357
transform 1 0 6074 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_270
timestamp 1717294357
transform 1 0 5285 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_271
timestamp 1717294357
transform 1 0 5126 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_272
timestamp 1717294357
transform 1 0 7022 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_273
timestamp 1717294357
transform 1 0 7338 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_274
timestamp 1717294357
transform 1 0 6390 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_275
timestamp 1717294357
transform 1 0 6706 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_276
timestamp 1717294357
transform 1 0 5442 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_277
timestamp 1717294357
transform 1 0 6074 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_278
timestamp 1717294357
transform 1 0 5758 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_279
timestamp 1717294357
transform 1 0 5126 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_280
timestamp 1717294357
transform 1 0 7181 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_281
timestamp 1717294357
transform 1 0 7497 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_282
timestamp 1717294357
transform 1 0 6233 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_283
timestamp 1717294357
transform 1 0 6549 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_284
timestamp 1717294357
transform 1 0 6865 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_285
timestamp 1717294357
transform 1 0 5601 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_286
timestamp 1717294357
transform 1 0 5917 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_287
timestamp 1717294357
transform 1 0 5285 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_288
timestamp 1717294357
transform 1 0 7022 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_289
timestamp 1717294357
transform 1 0 7338 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_290
timestamp 1717294357
transform 1 0 7181 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_291
timestamp 1717294357
transform 1 0 7497 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_292
timestamp 1717294357
transform 1 0 6390 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_293
timestamp 1717294357
transform 1 0 6233 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_294
timestamp 1717294357
transform 1 0 6706 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_295
timestamp 1717294357
transform 1 0 6549 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_296
timestamp 1717294357
transform 1 0 6865 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_297
timestamp 1717294357
transform 1 0 5442 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_298
timestamp 1717294357
transform 1 0 6074 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_299
timestamp 1717294357
transform 1 0 5758 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_300
timestamp 1717294357
transform 1 0 5601 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_301
timestamp 1717294357
transform 1 0 5917 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_302
timestamp 1717294357
transform 1 0 5126 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_303
timestamp 1717294357
transform 1 0 5285 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_304
timestamp 1717294357
transform 1 0 7022 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_305
timestamp 1717294357
transform 1 0 7338 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_306
timestamp 1717294357
transform 1 0 6390 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_307
timestamp 1717294357
transform 1 0 6706 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_308
timestamp 1717294357
transform 1 0 5442 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_309
timestamp 1717294357
transform 1 0 6074 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_310
timestamp 1717294357
transform 1 0 5758 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_311
timestamp 1717294357
transform 1 0 5126 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_312
timestamp 1717294357
transform 1 0 7181 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_313
timestamp 1717294357
transform 1 0 7497 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_314
timestamp 1717294357
transform 1 0 6233 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_315
timestamp 1717294357
transform 1 0 6549 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_316
timestamp 1717294357
transform 1 0 6865 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_317
timestamp 1717294357
transform 1 0 5601 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_318
timestamp 1717294357
transform 1 0 5917 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_319
timestamp 1717294357
transform 1 0 5285 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_320
timestamp 1717294357
transform 1 0 7181 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_321
timestamp 1717294357
transform 1 0 7497 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_322
timestamp 1717294357
transform 1 0 7022 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_323
timestamp 1717294357
transform 1 0 7338 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_324
timestamp 1717294357
transform 1 0 6233 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_325
timestamp 1717294357
transform 1 0 6390 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_326
timestamp 1717294357
transform 1 0 6549 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_327
timestamp 1717294357
transform 1 0 6865 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_328
timestamp 1717294357
transform 1 0 6706 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_329
timestamp 1717294357
transform 1 0 5601 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_330
timestamp 1717294357
transform 1 0 5917 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_331
timestamp 1717294357
transform 1 0 5442 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_332
timestamp 1717294357
transform 1 0 5758 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_333
timestamp 1717294357
transform 1 0 6074 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_334
timestamp 1717294357
transform 1 0 5285 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_335
timestamp 1717294357
transform 1 0 5126 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_336
timestamp 1717294357
transform 1 0 4494 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_337
timestamp 1717294357
transform 1 0 4810 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_338
timestamp 1717294357
transform 1 0 4653 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_339
timestamp 1717294357
transform 1 0 4337 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_340
timestamp 1717294357
transform 1 0 5442 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_341
timestamp 1717294357
transform 1 0 5758 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_342
timestamp 1717294357
transform 1 0 6074 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_343
timestamp 1717294357
transform 1 0 5126 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_344
timestamp 1717294357
transform 1 0 5601 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_345
timestamp 1717294357
transform 1 0 5917 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_346
timestamp 1717294357
transform 1 0 4969 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_347
timestamp 1717294357
transform 1 0 5285 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_348
timestamp 1717294357
transform 1 0 7022 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_349
timestamp 1717294357
transform 1 0 7338 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_350
timestamp 1717294357
transform 1 0 6390 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_351
timestamp 1717294357
transform 1 0 6706 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_352
timestamp 1717294357
transform 1 0 7181 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_353
timestamp 1717294357
transform 1 0 6233 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_354
timestamp 1717294357
transform 1 0 6865 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_355
timestamp 1717294357
transform 1 0 6549 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_356
timestamp 1717294357
transform 1 0 7497 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_357
timestamp 1717294357
transform 1 0 4494 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_358
timestamp 1717294357
transform 1 0 4810 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_359
timestamp 1717294357
transform 1 0 4653 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_360
timestamp 1717294357
transform 1 0 4337 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_361
timestamp 1717294357
transform 1 0 5442 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_362
timestamp 1717294357
transform 1 0 5758 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_363
timestamp 1717294357
transform 1 0 6074 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_364
timestamp 1717294357
transform 1 0 5126 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_365
timestamp 1717294357
transform 1 0 5601 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_366
timestamp 1717294357
transform 1 0 5917 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_367
timestamp 1717294357
transform 1 0 4969 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_368
timestamp 1717294357
transform 1 0 5285 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_369
timestamp 1717294357
transform 1 0 7022 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_370
timestamp 1717294357
transform 1 0 7338 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_371
timestamp 1717294357
transform 1 0 6390 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_372
timestamp 1717294357
transform 1 0 6706 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_373
timestamp 1717294357
transform 1 0 7181 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_374
timestamp 1717294357
transform 1 0 6233 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_375
timestamp 1717294357
transform 1 0 6865 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_376
timestamp 1717294357
transform 1 0 6549 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_377
timestamp 1717294357
transform 1 0 7497 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_378
timestamp 1717294357
transform 1 0 4653 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_379
timestamp 1717294357
transform 1 0 4494 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_380
timestamp 1717294357
transform 1 0 4810 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_381
timestamp 1717294357
transform 1 0 4337 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_382
timestamp 1717294357
transform 1 0 5601 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_383
timestamp 1717294357
transform 1 0 5917 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_384
timestamp 1717294357
transform 1 0 5442 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_385
timestamp 1717294357
transform 1 0 5758 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_386
timestamp 1717294357
transform 1 0 6074 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_387
timestamp 1717294357
transform 1 0 4969 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_388
timestamp 1717294357
transform 1 0 5285 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_389
timestamp 1717294357
transform 1 0 5126 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_390
timestamp 1717294357
transform 1 0 7181 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_391
timestamp 1717294357
transform 1 0 7022 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_392
timestamp 1717294357
transform 1 0 7338 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_393
timestamp 1717294357
transform 1 0 6233 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_394
timestamp 1717294357
transform 1 0 6390 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_395
timestamp 1717294357
transform 1 0 6865 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_396
timestamp 1717294357
transform 1 0 6549 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_397
timestamp 1717294357
transform 1 0 6706 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_398
timestamp 1717294357
transform 1 0 7497 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_399
timestamp 1717294357
transform 1 0 4653 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_400
timestamp 1717294357
transform 1 0 4337 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_401
timestamp 1717294357
transform 1 0 5917 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_402
timestamp 1717294357
transform 1 0 5601 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_403
timestamp 1717294357
transform 1 0 5285 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_404
timestamp 1717294357
transform 1 0 4969 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_405
timestamp 1717294357
transform 1 0 7181 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_406
timestamp 1717294357
transform 1 0 6233 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_407
timestamp 1717294357
transform 1 0 6549 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_408
timestamp 1717294357
transform 1 0 6865 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_409
timestamp 1717294357
transform 1 0 7497 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_410
timestamp 1717294357
transform 1 0 6390 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_411
timestamp 1717294357
transform 1 0 6706 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_412
timestamp 1717294357
transform 1 0 5758 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_413
timestamp 1717294357
transform 1 0 6074 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_414
timestamp 1717294357
transform 1 0 5442 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_415
timestamp 1717294357
transform 1 0 5126 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_416
timestamp 1717294357
transform 1 0 4810 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_417
timestamp 1717294357
transform 1 0 4494 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_418
timestamp 1717294357
transform 1 0 3890 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_419
timestamp 1717294357
transform 1 0 3574 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_420
timestamp 1717294357
transform 1 0 9206 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_421
timestamp 1717294357
transform 1 0 9522 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_422
timestamp 1717294357
transform 1 0 8890 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_423
timestamp 1717294357
transform 1 0 7942 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_424
timestamp 1717294357
transform 1 0 8574 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_425
timestamp 1717294357
transform 1 0 8258 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_426
timestamp 1717294357
transform 1 0 9681 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_427
timestamp 1717294357
transform 1 0 9365 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_428
timestamp 1717294357
transform 1 0 9049 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_429
timestamp 1717294357
transform 1 0 8733 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_430
timestamp 1717294357
transform 1 0 8101 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_431
timestamp 1717294357
transform 1 0 8417 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_432
timestamp 1717294357
transform 1 0 7785 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_433
timestamp 1717294357
transform 1 0 10470 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_434
timestamp 1717294357
transform 1 0 10786 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_435
timestamp 1717294357
transform 1 0 9838 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_436
timestamp 1717294357
transform 1 0 10154 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_437
timestamp 1717294357
transform 1 0 10629 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_438
timestamp 1717294357
transform 1 0 10945 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_439
timestamp 1717294357
transform 1 0 10313 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_440
timestamp 1717294357
transform 1 0 9997 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_441
timestamp 1717294357
transform 1 0 7785 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_442
timestamp 1717294357
transform 1 0 8101 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_443
timestamp 1717294357
transform 1 0 7942 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_444
timestamp 1717294357
transform 1 0 7785 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_445
timestamp 1717294357
transform 1 0 8101 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_446
timestamp 1717294357
transform 1 0 7942 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_447
timestamp 1717294357
transform 1 0 7785 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_448
timestamp 1717294357
transform 1 0 8101 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_449
timestamp 1717294357
transform 1 0 7942 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_450
timestamp 1717294357
transform 1 0 7785 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_451
timestamp 1717294357
transform 1 0 8101 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_452
timestamp 1717294357
transform 1 0 7942 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_453
timestamp 1717294357
transform 1 0 7785 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_454
timestamp 1717294357
transform 1 0 8101 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_455
timestamp 1717294357
transform 1 0 7942 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_456
timestamp 1717294357
transform 1 0 10629 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_457
timestamp 1717294357
transform 1 0 10945 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_458
timestamp 1717294357
transform 1 0 10470 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_459
timestamp 1717294357
transform 1 0 10786 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_460
timestamp 1717294357
transform 1 0 9997 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_461
timestamp 1717294357
transform 1 0 9681 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_462
timestamp 1717294357
transform 1 0 10313 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_463
timestamp 1717294357
transform 1 0 9838 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_464
timestamp 1717294357
transform 1 0 10154 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_465
timestamp 1717294357
transform 1 0 9365 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_466
timestamp 1717294357
transform 1 0 9522 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_467
timestamp 1717294357
transform 1 0 9206 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_468
timestamp 1717294357
transform 1 0 9049 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_469
timestamp 1717294357
transform 1 0 8890 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_470
timestamp 1717294357
transform 1 0 8733 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_471
timestamp 1717294357
transform 1 0 8417 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_472
timestamp 1717294357
transform 1 0 8258 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_473
timestamp 1717294357
transform 1 0 8574 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_474
timestamp 1717294357
transform 1 0 10470 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_475
timestamp 1717294357
transform 1 0 10786 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_476
timestamp 1717294357
transform 1 0 9838 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_477
timestamp 1717294357
transform 1 0 10154 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_478
timestamp 1717294357
transform 1 0 9522 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_479
timestamp 1717294357
transform 1 0 9206 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_480
timestamp 1717294357
transform 1 0 8890 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_481
timestamp 1717294357
transform 1 0 8258 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_482
timestamp 1717294357
transform 1 0 8574 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_483
timestamp 1717294357
transform 1 0 10629 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_484
timestamp 1717294357
transform 1 0 10945 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_485
timestamp 1717294357
transform 1 0 9681 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_486
timestamp 1717294357
transform 1 0 9997 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_487
timestamp 1717294357
transform 1 0 10313 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_488
timestamp 1717294357
transform 1 0 9365 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_489
timestamp 1717294357
transform 1 0 9049 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_490
timestamp 1717294357
transform 1 0 8733 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_491
timestamp 1717294357
transform 1 0 8417 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_492
timestamp 1717294357
transform 1 0 10470 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_493
timestamp 1717294357
transform 1 0 10786 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_494
timestamp 1717294357
transform 1 0 10629 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_495
timestamp 1717294357
transform 1 0 10945 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_496
timestamp 1717294357
transform 1 0 9838 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_497
timestamp 1717294357
transform 1 0 9681 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_498
timestamp 1717294357
transform 1 0 10154 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_499
timestamp 1717294357
transform 1 0 9997 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_500
timestamp 1717294357
transform 1 0 10313 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_501
timestamp 1717294357
transform 1 0 9522 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_502
timestamp 1717294357
transform 1 0 9206 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_503
timestamp 1717294357
transform 1 0 9365 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_504
timestamp 1717294357
transform 1 0 8890 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_505
timestamp 1717294357
transform 1 0 9049 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_506
timestamp 1717294357
transform 1 0 8733 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_507
timestamp 1717294357
transform 1 0 8258 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_508
timestamp 1717294357
transform 1 0 8574 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_509
timestamp 1717294357
transform 1 0 8417 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_510
timestamp 1717294357
transform 1 0 10470 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_511
timestamp 1717294357
transform 1 0 10786 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_512
timestamp 1717294357
transform 1 0 9838 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_513
timestamp 1717294357
transform 1 0 10154 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_514
timestamp 1717294357
transform 1 0 9522 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_515
timestamp 1717294357
transform 1 0 9206 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_516
timestamp 1717294357
transform 1 0 8890 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_517
timestamp 1717294357
transform 1 0 8574 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_518
timestamp 1717294357
transform 1 0 8258 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_519
timestamp 1717294357
transform 1 0 10629 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_520
timestamp 1717294357
transform 1 0 10945 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_521
timestamp 1717294357
transform 1 0 9681 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_522
timestamp 1717294357
transform 1 0 9997 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_523
timestamp 1717294357
transform 1 0 10313 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_524
timestamp 1717294357
transform 1 0 9365 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_525
timestamp 1717294357
transform 1 0 9049 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_526
timestamp 1717294357
transform 1 0 8733 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_527
timestamp 1717294357
transform 1 0 8417 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_528
timestamp 1717294357
transform 1 0 10629 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_529
timestamp 1717294357
transform 1 0 10945 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_530
timestamp 1717294357
transform 1 0 10470 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_531
timestamp 1717294357
transform 1 0 10786 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_532
timestamp 1717294357
transform 1 0 9681 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_533
timestamp 1717294357
transform 1 0 9838 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_534
timestamp 1717294357
transform 1 0 9997 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_535
timestamp 1717294357
transform 1 0 10313 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_536
timestamp 1717294357
transform 1 0 10154 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_537
timestamp 1717294357
transform 1 0 9365 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_538
timestamp 1717294357
transform 1 0 9206 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_539
timestamp 1717294357
transform 1 0 9522 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_540
timestamp 1717294357
transform 1 0 9049 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_541
timestamp 1717294357
transform 1 0 8890 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_542
timestamp 1717294357
transform 1 0 8733 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_543
timestamp 1717294357
transform 1 0 8417 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_544
timestamp 1717294357
transform 1 0 8258 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_545
timestamp 1717294357
transform 1 0 8574 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_546
timestamp 1717294357
transform 1 0 7942 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_547
timestamp 1717294357
transform 1 0 7785 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_548
timestamp 1717294357
transform 1 0 7942 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_549
timestamp 1717294357
transform 1 0 7785 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_550
timestamp 1717294357
transform 1 0 7942 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_551
timestamp 1717294357
transform 1 0 7785 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_552
timestamp 1717294357
transform 1 0 7785 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_553
timestamp 1717294357
transform 1 0 10629 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_554
timestamp 1717294357
transform 1 0 10945 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_555
timestamp 1717294357
transform 1 0 9681 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_556
timestamp 1717294357
transform 1 0 9997 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_557
timestamp 1717294357
transform 1 0 10313 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_558
timestamp 1717294357
transform 1 0 9365 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_559
timestamp 1717294357
transform 1 0 9049 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_560
timestamp 1717294357
transform 1 0 8733 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_561
timestamp 1717294357
transform 1 0 8101 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_562
timestamp 1717294357
transform 1 0 8417 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_563
timestamp 1717294357
transform 1 0 10945 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_564
timestamp 1717294357
transform 1 0 10629 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_565
timestamp 1717294357
transform 1 0 10470 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_566
timestamp 1717294357
transform 1 0 10786 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_567
timestamp 1717294357
transform 1 0 9997 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_568
timestamp 1717294357
transform 1 0 9681 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_569
timestamp 1717294357
transform 1 0 10313 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_570
timestamp 1717294357
transform 1 0 9838 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_571
timestamp 1717294357
transform 1 0 10154 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_572
timestamp 1717294357
transform 1 0 9365 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_573
timestamp 1717294357
transform 1 0 9522 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_574
timestamp 1717294357
transform 1 0 9206 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_575
timestamp 1717294357
transform 1 0 9049 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_576
timestamp 1717294357
transform 1 0 8890 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_577
timestamp 1717294357
transform 1 0 8733 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_578
timestamp 1717294357
transform 1 0 8101 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_579
timestamp 1717294357
transform 1 0 8417 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_580
timestamp 1717294357
transform 1 0 8258 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_581
timestamp 1717294357
transform 1 0 8574 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_582
timestamp 1717294357
transform 1 0 10470 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_583
timestamp 1717294357
transform 1 0 10786 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_584
timestamp 1717294357
transform 1 0 9838 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_585
timestamp 1717294357
transform 1 0 10154 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_586
timestamp 1717294357
transform 1 0 9522 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_587
timestamp 1717294357
transform 1 0 9206 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_588
timestamp 1717294357
transform 1 0 8890 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_589
timestamp 1717294357
transform 1 0 8258 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_590
timestamp 1717294357
transform 1 0 8574 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_591
timestamp 1717294357
transform 1 0 10470 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_592
timestamp 1717294357
transform 1 0 10786 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_593
timestamp 1717294357
transform 1 0 10945 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_594
timestamp 1717294357
transform 1 0 10629 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_595
timestamp 1717294357
transform 1 0 9838 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_596
timestamp 1717294357
transform 1 0 10154 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_597
timestamp 1717294357
transform 1 0 9997 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_598
timestamp 1717294357
transform 1 0 9681 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_599
timestamp 1717294357
transform 1 0 10313 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_600
timestamp 1717294357
transform 1 0 9522 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_601
timestamp 1717294357
transform 1 0 9206 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_602
timestamp 1717294357
transform 1 0 9365 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_603
timestamp 1717294357
transform 1 0 8890 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_604
timestamp 1717294357
transform 1 0 9049 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_605
timestamp 1717294357
transform 1 0 8733 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_606
timestamp 1717294357
transform 1 0 8258 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_607
timestamp 1717294357
transform 1 0 8574 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_608
timestamp 1717294357
transform 1 0 8101 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_609
timestamp 1717294357
transform 1 0 8417 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_610
timestamp 1717294357
transform 1 0 10629 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_611
timestamp 1717294357
transform 1 0 10945 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_612
timestamp 1717294357
transform 1 0 9997 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_613
timestamp 1717294357
transform 1 0 9681 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_614
timestamp 1717294357
transform 1 0 10313 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_615
timestamp 1717294357
transform 1 0 9365 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_616
timestamp 1717294357
transform 1 0 9049 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_617
timestamp 1717294357
transform 1 0 8733 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_618
timestamp 1717294357
transform 1 0 8101 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_619
timestamp 1717294357
transform 1 0 8417 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_620
timestamp 1717294357
transform 1 0 7942 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_621
timestamp 1717294357
transform 1 0 10470 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_622
timestamp 1717294357
transform 1 0 10786 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_623
timestamp 1717294357
transform 1 0 9838 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_624
timestamp 1717294357
transform 1 0 10154 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_625
timestamp 1717294357
transform 1 0 9206 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_626
timestamp 1717294357
transform 1 0 9522 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_627
timestamp 1717294357
transform 1 0 12338 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_628
timestamp 1717294357
transform 1 0 12022 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_629
timestamp 1717294357
transform 1 0 11706 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_630
timestamp 1717294357
transform 1 0 12654 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_631
timestamp 1717294357
transform 1 0 12970 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_632
timestamp 1717294357
transform 1 0 12338 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_633
timestamp 1717294357
transform 1 0 11390 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_634
timestamp 1717294357
transform 1 0 12022 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_635
timestamp 1717294357
transform 1 0 11706 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_636
timestamp 1717294357
transform 1 0 13129 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_637
timestamp 1717294357
transform 1 0 12813 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_638
timestamp 1717294357
transform 1 0 12497 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_639
timestamp 1717294357
transform 1 0 12181 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_640
timestamp 1717294357
transform 1 0 11549 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_641
timestamp 1717294357
transform 1 0 11865 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_642
timestamp 1717294357
transform 1 0 11233 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_643
timestamp 1717294357
transform 1 0 13918 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_644
timestamp 1717294357
transform 1 0 14234 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_645
timestamp 1717294357
transform 1 0 13286 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_646
timestamp 1717294357
transform 1 0 13602 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_647
timestamp 1717294357
transform 1 0 14077 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_648
timestamp 1717294357
transform 1 0 14393 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_649
timestamp 1717294357
transform 1 0 13761 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_650
timestamp 1717294357
transform 1 0 13445 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_651
timestamp 1717294357
transform 1 0 11233 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_652
timestamp 1717294357
transform 1 0 11233 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_653
timestamp 1717294357
transform 1 0 11233 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_654
timestamp 1717294357
transform 1 0 11233 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_655
timestamp 1717294357
transform 1 0 11233 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_656
timestamp 1717294357
transform 1 0 14077 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_657
timestamp 1717294357
transform 1 0 14393 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_658
timestamp 1717294357
transform 1 0 13918 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_659
timestamp 1717294357
transform 1 0 14234 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_660
timestamp 1717294357
transform 1 0 13129 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_661
timestamp 1717294357
transform 1 0 13445 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_662
timestamp 1717294357
transform 1 0 13761 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_663
timestamp 1717294357
transform 1 0 13286 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_664
timestamp 1717294357
transform 1 0 13602 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_665
timestamp 1717294357
transform 1 0 12813 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_666
timestamp 1717294357
transform 1 0 12970 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_667
timestamp 1717294357
transform 1 0 12654 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_668
timestamp 1717294357
transform 1 0 12497 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_669
timestamp 1717294357
transform 1 0 12338 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_670
timestamp 1717294357
transform 1 0 12181 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_671
timestamp 1717294357
transform 1 0 11549 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_672
timestamp 1717294357
transform 1 0 11865 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_673
timestamp 1717294357
transform 1 0 11390 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_674
timestamp 1717294357
transform 1 0 11706 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_675
timestamp 1717294357
transform 1 0 12022 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_676
timestamp 1717294357
transform 1 0 13918 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_677
timestamp 1717294357
transform 1 0 14234 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_678
timestamp 1717294357
transform 1 0 13286 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_679
timestamp 1717294357
transform 1 0 13602 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_680
timestamp 1717294357
transform 1 0 12970 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_681
timestamp 1717294357
transform 1 0 12654 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_682
timestamp 1717294357
transform 1 0 12338 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_683
timestamp 1717294357
transform 1 0 11706 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_684
timestamp 1717294357
transform 1 0 12022 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_685
timestamp 1717294357
transform 1 0 11390 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_686
timestamp 1717294357
transform 1 0 14077 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_687
timestamp 1717294357
transform 1 0 14393 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_688
timestamp 1717294357
transform 1 0 13129 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_689
timestamp 1717294357
transform 1 0 13445 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_690
timestamp 1717294357
transform 1 0 13761 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_691
timestamp 1717294357
transform 1 0 12813 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_692
timestamp 1717294357
transform 1 0 12497 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_693
timestamp 1717294357
transform 1 0 12181 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_694
timestamp 1717294357
transform 1 0 11865 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_695
timestamp 1717294357
transform 1 0 11549 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_696
timestamp 1717294357
transform 1 0 13918 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_697
timestamp 1717294357
transform 1 0 14234 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_698
timestamp 1717294357
transform 1 0 14077 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_699
timestamp 1717294357
transform 1 0 14393 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_700
timestamp 1717294357
transform 1 0 13129 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_701
timestamp 1717294357
transform 1 0 13286 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_702
timestamp 1717294357
transform 1 0 13602 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_703
timestamp 1717294357
transform 1 0 13445 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_704
timestamp 1717294357
transform 1 0 13761 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_705
timestamp 1717294357
transform 1 0 12970 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_706
timestamp 1717294357
transform 1 0 12654 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_707
timestamp 1717294357
transform 1 0 12813 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_708
timestamp 1717294357
transform 1 0 12338 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_709
timestamp 1717294357
transform 1 0 12497 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_710
timestamp 1717294357
transform 1 0 12181 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_711
timestamp 1717294357
transform 1 0 11706 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_712
timestamp 1717294357
transform 1 0 12022 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_713
timestamp 1717294357
transform 1 0 11390 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_714
timestamp 1717294357
transform 1 0 11865 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_715
timestamp 1717294357
transform 1 0 11549 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_716
timestamp 1717294357
transform 1 0 13918 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_717
timestamp 1717294357
transform 1 0 14234 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_718
timestamp 1717294357
transform 1 0 13286 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_719
timestamp 1717294357
transform 1 0 13602 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_720
timestamp 1717294357
transform 1 0 12970 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_721
timestamp 1717294357
transform 1 0 12654 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_722
timestamp 1717294357
transform 1 0 12338 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_723
timestamp 1717294357
transform 1 0 12022 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_724
timestamp 1717294357
transform 1 0 11706 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_725
timestamp 1717294357
transform 1 0 11390 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_726
timestamp 1717294357
transform 1 0 14077 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_727
timestamp 1717294357
transform 1 0 14393 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_728
timestamp 1717294357
transform 1 0 13129 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_729
timestamp 1717294357
transform 1 0 13445 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_730
timestamp 1717294357
transform 1 0 13761 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_731
timestamp 1717294357
transform 1 0 12813 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_732
timestamp 1717294357
transform 1 0 12497 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_733
timestamp 1717294357
transform 1 0 12181 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_734
timestamp 1717294357
transform 1 0 11549 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_735
timestamp 1717294357
transform 1 0 11865 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_736
timestamp 1717294357
transform 1 0 14077 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_737
timestamp 1717294357
transform 1 0 14393 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_738
timestamp 1717294357
transform 1 0 13918 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_739
timestamp 1717294357
transform 1 0 14234 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_740
timestamp 1717294357
transform 1 0 13129 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_741
timestamp 1717294357
transform 1 0 13286 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_742
timestamp 1717294357
transform 1 0 13445 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_743
timestamp 1717294357
transform 1 0 13761 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_744
timestamp 1717294357
transform 1 0 13602 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_745
timestamp 1717294357
transform 1 0 12813 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_746
timestamp 1717294357
transform 1 0 12654 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_747
timestamp 1717294357
transform 1 0 12970 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_748
timestamp 1717294357
transform 1 0 12497 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_749
timestamp 1717294357
transform 1 0 12338 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_750
timestamp 1717294357
transform 1 0 12181 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_751
timestamp 1717294357
transform 1 0 11549 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_752
timestamp 1717294357
transform 1 0 11865 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_753
timestamp 1717294357
transform 1 0 11390 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_754
timestamp 1717294357
transform 1 0 11706 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_755
timestamp 1717294357
transform 1 0 12022 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_756
timestamp 1717294357
transform 1 0 11549 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_757
timestamp 1717294357
transform 1 0 11233 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_758
timestamp 1717294357
transform 1 0 12181 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_759
timestamp 1717294357
transform 1 0 11865 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_760
timestamp 1717294357
transform 1 0 11390 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_761
timestamp 1717294357
transform 1 0 11706 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_762
timestamp 1717294357
transform 1 0 12022 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_763
timestamp 1717294357
transform 1 0 12338 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_764
timestamp 1717294357
transform 1 0 11549 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_765
timestamp 1717294357
transform 1 0 11233 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_766
timestamp 1717294357
transform 1 0 12181 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_767
timestamp 1717294357
transform 1 0 11865 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_768
timestamp 1717294357
transform 1 0 11390 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_769
timestamp 1717294357
transform 1 0 11706 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_770
timestamp 1717294357
transform 1 0 12022 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_771
timestamp 1717294357
transform 1 0 12338 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_772
timestamp 1717294357
transform 1 0 11549 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_773
timestamp 1717294357
transform 1 0 11233 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_774
timestamp 1717294357
transform 1 0 12181 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_775
timestamp 1717294357
transform 1 0 11865 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_776
timestamp 1717294357
transform 1 0 11390 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_777
timestamp 1717294357
transform 1 0 11706 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_778
timestamp 1717294357
transform 1 0 12022 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_779
timestamp 1717294357
transform 1 0 12338 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_780
timestamp 1717294357
transform 1 0 11549 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_781
timestamp 1717294357
transform 1 0 11233 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_782
timestamp 1717294357
transform 1 0 12181 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_783
timestamp 1717294357
transform 1 0 11865 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_784
timestamp 1717294357
transform 1 0 14077 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_785
timestamp 1717294357
transform 1 0 14393 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_786
timestamp 1717294357
transform 1 0 13129 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_787
timestamp 1717294357
transform 1 0 13445 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_788
timestamp 1717294357
transform 1 0 13761 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_789
timestamp 1717294357
transform 1 0 12813 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_790
timestamp 1717294357
transform 1 0 12497 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_791
timestamp 1717294357
transform 1 0 14393 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_792
timestamp 1717294357
transform 1 0 14077 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_793
timestamp 1717294357
transform 1 0 13918 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_794
timestamp 1717294357
transform 1 0 14234 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_795
timestamp 1717294357
transform 1 0 13129 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_796
timestamp 1717294357
transform 1 0 13445 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_797
timestamp 1717294357
transform 1 0 13761 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_798
timestamp 1717294357
transform 1 0 13286 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_799
timestamp 1717294357
transform 1 0 13602 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_800
timestamp 1717294357
transform 1 0 12813 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_801
timestamp 1717294357
transform 1 0 12970 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_802
timestamp 1717294357
transform 1 0 12654 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_803
timestamp 1717294357
transform 1 0 12497 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_804
timestamp 1717294357
transform 1 0 13918 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_805
timestamp 1717294357
transform 1 0 14234 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_806
timestamp 1717294357
transform 1 0 13286 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_807
timestamp 1717294357
transform 1 0 13602 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_808
timestamp 1717294357
transform 1 0 12970 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_809
timestamp 1717294357
transform 1 0 12654 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_810
timestamp 1717294357
transform 1 0 13918 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_811
timestamp 1717294357
transform 1 0 14234 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_812
timestamp 1717294357
transform 1 0 14393 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_813
timestamp 1717294357
transform 1 0 14077 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_814
timestamp 1717294357
transform 1 0 13286 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_815
timestamp 1717294357
transform 1 0 13602 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_816
timestamp 1717294357
transform 1 0 13129 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_817
timestamp 1717294357
transform 1 0 13445 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_818
timestamp 1717294357
transform 1 0 13761 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_819
timestamp 1717294357
transform 1 0 12970 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_820
timestamp 1717294357
transform 1 0 12654 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_821
timestamp 1717294357
transform 1 0 12813 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_822
timestamp 1717294357
transform 1 0 12497 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_823
timestamp 1717294357
transform 1 0 14077 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_824
timestamp 1717294357
transform 1 0 14393 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_825
timestamp 1717294357
transform 1 0 13129 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_826
timestamp 1717294357
transform 1 0 13445 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_827
timestamp 1717294357
transform 1 0 13761 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_828
timestamp 1717294357
transform 1 0 12813 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_829
timestamp 1717294357
transform 1 0 12497 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_830
timestamp 1717294357
transform 1 0 11390 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_831
timestamp 1717294357
transform 1 0 8890 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_832
timestamp 1717294357
transform 1 0 8574 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_833
timestamp 1717294357
transform 1 0 8258 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_834
timestamp 1717294357
transform 1 0 13918 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_835
timestamp 1717294357
transform 1 0 14234 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_836
timestamp 1717294357
transform 1 0 13286 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_837
timestamp 1717294357
transform 1 0 13602 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_838
timestamp 1717294357
transform 1 0 16102 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_839
timestamp 1717294357
transform 1 0 16418 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_840
timestamp 1717294357
transform 1 0 16102 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_841
timestamp 1717294357
transform 1 0 16418 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_842
timestamp 1717294357
transform 1 0 15786 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_843
timestamp 1717294357
transform 1 0 14838 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_844
timestamp 1717294357
transform 1 0 15470 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_845
timestamp 1717294357
transform 1 0 15154 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_846
timestamp 1717294357
transform 1 0 16261 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_847
timestamp 1717294357
transform 1 0 15945 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_848
timestamp 1717294357
transform 1 0 15629 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_849
timestamp 1717294357
transform 1 0 14997 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_850
timestamp 1717294357
transform 1 0 15313 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_851
timestamp 1717294357
transform 1 0 14681 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_852
timestamp 1717294357
transform 1 0 17366 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_853
timestamp 1717294357
transform 1 0 17682 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_854
timestamp 1717294357
transform 1 0 16734 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_855
timestamp 1717294357
transform 1 0 17050 0 1 496
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_856
timestamp 1717294357
transform 1 0 17525 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_857
timestamp 1717294357
transform 1 0 17841 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_858
timestamp 1717294357
transform 1 0 16577 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_859
timestamp 1717294357
transform 1 0 17209 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_860
timestamp 1717294357
transform 1 0 16893 0 1 -4
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_861
timestamp 1717294357
transform 1 0 17525 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_862
timestamp 1717294357
transform 1 0 17366 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_863
timestamp 1717294357
transform 1 0 16577 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_864
timestamp 1717294357
transform 1 0 16893 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_865
timestamp 1717294357
transform 1 0 17209 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_866
timestamp 1717294357
transform 1 0 16734 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_867
timestamp 1717294357
transform 1 0 17050 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_868
timestamp 1717294357
transform 1 0 16261 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_869
timestamp 1717294357
transform 1 0 16418 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_870
timestamp 1717294357
transform 1 0 16102 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_871
timestamp 1717294357
transform 1 0 15945 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_872
timestamp 1717294357
transform 1 0 15786 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_873
timestamp 1717294357
transform 1 0 15629 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_874
timestamp 1717294357
transform 1 0 14997 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_875
timestamp 1717294357
transform 1 0 15313 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_876
timestamp 1717294357
transform 1 0 14838 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_877
timestamp 1717294357
transform 1 0 15154 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_878
timestamp 1717294357
transform 1 0 15470 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_879
timestamp 1717294357
transform 1 0 14681 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_880
timestamp 1717294357
transform 1 0 17366 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_881
timestamp 1717294357
transform 1 0 16734 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_882
timestamp 1717294357
transform 1 0 17050 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_883
timestamp 1717294357
transform 1 0 16418 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_884
timestamp 1717294357
transform 1 0 16102 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_885
timestamp 1717294357
transform 1 0 15786 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_886
timestamp 1717294357
transform 1 0 15154 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_887
timestamp 1717294357
transform 1 0 15470 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_888
timestamp 1717294357
transform 1 0 14838 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_889
timestamp 1717294357
transform 1 0 17525 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_890
timestamp 1717294357
transform 1 0 16577 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_891
timestamp 1717294357
transform 1 0 16893 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_892
timestamp 1717294357
transform 1 0 17209 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_893
timestamp 1717294357
transform 1 0 16261 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_894
timestamp 1717294357
transform 1 0 15945 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_895
timestamp 1717294357
transform 1 0 15629 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_896
timestamp 1717294357
transform 1 0 15313 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_897
timestamp 1717294357
transform 1 0 14997 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_898
timestamp 1717294357
transform 1 0 14681 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_899
timestamp 1717294357
transform 1 0 17366 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_900
timestamp 1717294357
transform 1 0 17525 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_901
timestamp 1717294357
transform 1 0 16577 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_902
timestamp 1717294357
transform 1 0 16734 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_903
timestamp 1717294357
transform 1 0 17050 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_904
timestamp 1717294357
transform 1 0 16893 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_905
timestamp 1717294357
transform 1 0 17209 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_906
timestamp 1717294357
transform 1 0 16418 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_907
timestamp 1717294357
transform 1 0 16102 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_908
timestamp 1717294357
transform 1 0 16261 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_909
timestamp 1717294357
transform 1 0 15786 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_910
timestamp 1717294357
transform 1 0 15945 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_911
timestamp 1717294357
transform 1 0 15629 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_912
timestamp 1717294357
transform 1 0 15154 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_913
timestamp 1717294357
transform 1 0 15470 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_914
timestamp 1717294357
transform 1 0 14838 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_915
timestamp 1717294357
transform 1 0 15313 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_916
timestamp 1717294357
transform 1 0 14997 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_917
timestamp 1717294357
transform 1 0 14681 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_918
timestamp 1717294357
transform 1 0 17366 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_919
timestamp 1717294357
transform 1 0 16734 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_920
timestamp 1717294357
transform 1 0 17050 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_921
timestamp 1717294357
transform 1 0 16418 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_922
timestamp 1717294357
transform 1 0 16102 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_923
timestamp 1717294357
transform 1 0 15786 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_924
timestamp 1717294357
transform 1 0 15470 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_925
timestamp 1717294357
transform 1 0 15154 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_926
timestamp 1717294357
transform 1 0 14838 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_927
timestamp 1717294357
transform 1 0 17525 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_928
timestamp 1717294357
transform 1 0 16577 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_929
timestamp 1717294357
transform 1 0 16893 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_930
timestamp 1717294357
transform 1 0 17209 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_931
timestamp 1717294357
transform 1 0 16261 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_932
timestamp 1717294357
transform 1 0 15945 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_933
timestamp 1717294357
transform 1 0 15629 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_934
timestamp 1717294357
transform 1 0 14997 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_935
timestamp 1717294357
transform 1 0 15313 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_936
timestamp 1717294357
transform 1 0 14681 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_937
timestamp 1717294357
transform 1 0 17525 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_938
timestamp 1717294357
transform 1 0 17366 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_939
timestamp 1717294357
transform 1 0 16577 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_940
timestamp 1717294357
transform 1 0 16734 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_941
timestamp 1717294357
transform 1 0 16893 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_942
timestamp 1717294357
transform 1 0 17209 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_943
timestamp 1717294357
transform 1 0 17050 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_944
timestamp 1717294357
transform 1 0 16261 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_945
timestamp 1717294357
transform 1 0 16102 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_946
timestamp 1717294357
transform 1 0 16418 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_947
timestamp 1717294357
transform 1 0 15945 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_948
timestamp 1717294357
transform 1 0 15786 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_949
timestamp 1717294357
transform 1 0 15629 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_950
timestamp 1717294357
transform 1 0 14997 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_951
timestamp 1717294357
transform 1 0 15313 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_952
timestamp 1717294357
transform 1 0 14838 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_953
timestamp 1717294357
transform 1 0 15154 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_954
timestamp 1717294357
transform 1 0 15470 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_955
timestamp 1717294357
transform 1 0 14681 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_956
timestamp 1717294357
transform 1 0 17682 0 1 6586
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_957
timestamp 1717294357
transform 1 0 17841 0 1 6086
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_958
timestamp 1717294357
transform 1 0 17682 0 1 5368
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_959
timestamp 1717294357
transform 1 0 17841 0 1 4868
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_960
timestamp 1717294357
transform 1 0 17682 0 1 4150
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_961
timestamp 1717294357
transform 1 0 17841 0 1 3650
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_962
timestamp 1717294357
transform 1 0 17682 0 1 2932
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_963
timestamp 1717294357
transform 1 0 17841 0 1 2432
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_964
timestamp 1717294357
transform 1 0 17682 0 1 1714
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_965
timestamp 1717294357
transform 1 0 17841 0 1 1214
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_966
timestamp 1717294357
transform 1 0 14681 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_967
timestamp 1717294357
transform 1 0 14997 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_968
timestamp 1717294357
transform 1 0 15313 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_969
timestamp 1717294357
transform 1 0 15945 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_970
timestamp 1717294357
transform 1 0 15629 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_971
timestamp 1717294357
transform 1 0 16577 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_972
timestamp 1717294357
transform 1 0 16261 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_973
timestamp 1717294357
transform 1 0 14838 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_974
timestamp 1717294357
transform 1 0 15154 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_975
timestamp 1717294357
transform 1 0 15470 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_976
timestamp 1717294357
transform 1 0 16102 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_977
timestamp 1717294357
transform 1 0 15786 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_978
timestamp 1717294357
transform 1 0 16418 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_979
timestamp 1717294357
transform 1 0 14681 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_980
timestamp 1717294357
transform 1 0 14997 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_981
timestamp 1717294357
transform 1 0 15313 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_982
timestamp 1717294357
transform 1 0 15945 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_983
timestamp 1717294357
transform 1 0 15629 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_984
timestamp 1717294357
transform 1 0 16577 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_985
timestamp 1717294357
transform 1 0 16261 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_986
timestamp 1717294357
transform 1 0 14838 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_987
timestamp 1717294357
transform 1 0 15154 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_988
timestamp 1717294357
transform 1 0 15470 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_989
timestamp 1717294357
transform 1 0 16102 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_990
timestamp 1717294357
transform 1 0 15786 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_991
timestamp 1717294357
transform 1 0 16418 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_992
timestamp 1717294357
transform 1 0 14681 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_993
timestamp 1717294357
transform 1 0 14997 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_994
timestamp 1717294357
transform 1 0 15313 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_995
timestamp 1717294357
transform 1 0 15945 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_996
timestamp 1717294357
transform 1 0 15629 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_997
timestamp 1717294357
transform 1 0 16577 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_998
timestamp 1717294357
transform 1 0 16261 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_999
timestamp 1717294357
transform 1 0 14838 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1000
timestamp 1717294357
transform 1 0 15154 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1001
timestamp 1717294357
transform 1 0 15470 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1002
timestamp 1717294357
transform 1 0 16102 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1003
timestamp 1717294357
transform 1 0 15786 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1004
timestamp 1717294357
transform 1 0 16418 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1005
timestamp 1717294357
transform 1 0 14681 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1006
timestamp 1717294357
transform 1 0 14997 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1007
timestamp 1717294357
transform 1 0 15313 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1008
timestamp 1717294357
transform 1 0 15945 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1009
timestamp 1717294357
transform 1 0 15629 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1010
timestamp 1717294357
transform 1 0 16577 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1011
timestamp 1717294357
transform 1 0 16261 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1012
timestamp 1717294357
transform 1 0 17525 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1013
timestamp 1717294357
transform 1 0 17841 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1014
timestamp 1717294357
transform 1 0 16893 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1015
timestamp 1717294357
transform 1 0 17209 0 1 10958
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1016
timestamp 1717294357
transform 1 0 17525 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1017
timestamp 1717294357
transform 1 0 17366 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1018
timestamp 1717294357
transform 1 0 17682 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1019
timestamp 1717294357
transform 1 0 17841 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1020
timestamp 1717294357
transform 1 0 16893 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1021
timestamp 1717294357
transform 1 0 17209 0 1 9740
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1022
timestamp 1717294357
transform 1 0 16734 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1023
timestamp 1717294357
transform 1 0 17050 0 1 10240
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1024
timestamp 1717294357
transform 1 0 17366 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1025
timestamp 1717294357
transform 1 0 17682 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1026
timestamp 1717294357
transform 1 0 16734 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1027
timestamp 1717294357
transform 1 0 17050 0 1 9022
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1028
timestamp 1717294357
transform 1 0 17366 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1029
timestamp 1717294357
transform 1 0 17682 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1030
timestamp 1717294357
transform 1 0 17525 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1031
timestamp 1717294357
transform 1 0 17841 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1032
timestamp 1717294357
transform 1 0 16734 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1033
timestamp 1717294357
transform 1 0 17050 0 1 7804
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1034
timestamp 1717294357
transform 1 0 16893 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1035
timestamp 1717294357
transform 1 0 17209 0 1 8522
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1036
timestamp 1717294357
transform 1 0 17525 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1037
timestamp 1717294357
transform 1 0 17841 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1038
timestamp 1717294357
transform 1 0 16893 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1039
timestamp 1717294357
transform 1 0 17209 0 1 7304
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1040
timestamp 1717294357
transform 1 0 15786 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1041
timestamp 1717294357
transform 1 0 15470 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1042
timestamp 1717294357
transform 1 0 15154 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1043
timestamp 1717294357
transform 1 0 14838 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1044
timestamp 1717294357
transform 1 0 12654 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1045
timestamp 1717294357
transform 1 0 12970 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1046
timestamp 1717294357
transform 1 0 17366 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1047
timestamp 1717294357
transform 1 0 17682 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1048
timestamp 1717294357
transform 1 0 16734 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1049
timestamp 1717294357
transform 1 0 17050 0 1 11458
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1050
timestamp 1717294357
transform 1 0 -2584 0 1 10654
box 9158 -5776 9224 -5362
use ldo_via_6cut  ldo_via_6cut_1051
timestamp 1717294357
transform 1 0 -4696 0 1 10645
box 9158 -5776 9224 -5362
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  sky130_fd_pr__pfet_g5v0d10v5_KLAZY6_0 paramcells
timestamp 1717294357
transform 1 0 5888 0 1 -6196
box -308 -397 308 397
use sky130_fd_sc_hvl__lsbuflv2hv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform -1 0 6586 0 -1 6296
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  x2
timestamp 1723858470
transform -1 0 8698 0 -1 6296
box -66 -43 2178 1671
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC1 paramcells
array 0 0 -1051 0 2 3379
timestamp 1717294357
transform -1 0 6647 0 1 -4177
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC3 paramcells
timestamp 1717294357
transform -1 0 5647 0 1 -9441
box -686 -540 686 540
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM46 paramcells
timestamp 1717294357
transform 1 0 5642 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__nfet_g5v0d10v5_69K6TN  XM48 paramcells
timestamp 1717294357
transform 1 0 9294 0 1 -8726
box -938 -358 938 358
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0  XM52 paramcells
timestamp 1717294357
transform 1 0 7902 0 1 -8240
box -288 -458 288 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0  XM53
timestamp 1717294357
transform 1 0 7456 0 1 -8240
box -288 -458 288 458
use sky130_fd_pr__nfet_g5v0d10v5_L9TFKV  XM54 paramcells
timestamp 1717294357
transform 1 0 5860 0 1 -8340
box -1128 -558 1128 558
use sky130_fd_pr__nfet_g5v0d10v5_69K6TN  XM55
timestamp 1717294357
transform 1 0 9294 0 1 -8140
box -938 -358 938 358
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM56
timestamp 1717294357
transform 1 0 7794 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM57
timestamp 1717294357
transform 1 0 8870 0 1 -7247
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM58
timestamp 1717294357
transform 1 0 6718 0 1 -7247
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM59
timestamp 1717294357
transform 1 0 11022 0 1 -7247
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM60
timestamp 1717294357
transform 1 0 9946 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__nfet_g5v0d10v5_YHRXVR  XM61 paramcells
array 0 4 3448 0 0 12478
timestamp 1717294357
transform 1 0 11659 0 1 156
box -1789 -6239 1789 6239
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM62
timestamp 1717294357
transform -1 0 18302 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM63
timestamp 1717294357
transform -1 0 19378 0 1 -7247
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM64
timestamp 1717294357
transform -1 0 16150 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM65
timestamp 1717294357
transform -1 0 17226 0 1 -7247
box -308 -397 308 397
use sky130_fd_pr__nfet_g5v0d10v5_A2FZRM  XM66 paramcells
array 0 3 2146 0 0 2388
timestamp 1717294357
transform 1 0 18252 0 1 -8972
box -1138 -1194 1138 1194
use sky130_fd_pr__nfet_g5v0d10v5_A2FZRM  XM67
timestamp 1717294357
transform 1 0 16106 0 1 -8972
box -1138 -1194 1138 1194
use sky130_fd_pr__pfet_g5v0d10v5_PC2PN5  XM68 paramcells
timestamp 1717294357
transform 1 0 14124 0 1 -7247
box -1258 -397 1258 397
use sky130_fd_pr__nfet_g5v0d10v5_A2FZRM  XM69
timestamp 1717294357
transform 1 0 13960 0 1 -8972
box -1138 -1194 1138 1194
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM70 paramcells
timestamp 1717294357
transform 1 0 27564 0 1 -7244
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_47NWVV  XM71 paramcells
timestamp 1717294357
transform 1 0 21406 0 1 -7247
box -458 -397 458 397
use sky130_fd_pr__pfet_g5v0d10v5_47NWVV  XM72
timestamp 1717294357
transform 1 0 20680 0 1 -7247
box -458 -397 458 397
use sky130_fd_pr__pfet_g5v0d10v5_47NWVV  XM73
timestamp 1717294357
transform 1 0 19954 0 1 -7247
box -458 -397 458 397
use sky130_fd_pr__nfet_g5v0d10v5_A2FZRM  XM74
timestamp 1717294357
transform 1 0 26836 0 1 -8972
box -1138 -1194 1138 1194
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM75
timestamp 1717294357
transform 1 0 7455 0 1 -9169
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6  XM76 paramcells
timestamp 1717294357
transform 1 0 5730 0 1 -9507
box -308 -547 308 547
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM77
timestamp 1717294357
transform 1 0 7901 0 1 -9169
box -288 -358 288 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM78
timestamp 1717294357
transform 1 0 7455 0 1 -9755
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_BWAZV5  XM79
timestamp 1717294357
transform 1 0 12098 0 1 -7247
box -958 -397 958 397
use sky130_fd_pr__nfet_g5v0d10v5_PXBJUB  XM80 paramcells
timestamp 1717294357
transform 1 0 11594 0 1 -8722
box -1228 -358 1228 358
use sky130_fd_pr__nfet_g5v0d10v5_PXBJUB  XM81
timestamp 1717294357
transform 1 0 11594 0 1 -8136
box -1228 -358 1228 358
use sky130_fd_pr__nfet_g5v0d10v5_PXBJUB  XM82
timestamp 1717294357
transform 1 0 11594 0 1 -9308
box -1228 -358 1228 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM83
timestamp 1717294357
transform 1 0 7901 0 1 -9755
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6  XM84
timestamp 1717294357
transform 1 0 6156 0 1 -9507
box -308 -547 308 547
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM85
timestamp 1717294357
transform 1 0 8915 0 1 -9609
box -288 -358 288 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM87
timestamp 1717294357
transform 1 0 9361 0 1 -9609
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM88
timestamp 1717294357
transform 1 0 6314 0 1 -6196
box -308 -397 308 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM89
timestamp 1717294357
transform 1 0 9807 0 1 -9609
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM90
timestamp 1717294357
transform 1 0 6740 0 1 -6196
box -308 -397 308 397
use sky130_fd_pr__res_xhigh_po_0p35_QZEXQH  XR4 paramcells
timestamp 1717294357
transform 0 1 6535 1 0 2264
box -1612 -1582 1612 1582
use sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H  XR5 paramcells
timestamp 1717294357
transform 0 1 6533 1 0 -2522
box -3106 -1582 3106 1582
use sky130_fd_pr__res_xhigh_po_0p35_743D3R  XR6 paramcells
timestamp 1717294357
transform 0 1 24580 -1 0 -7318
box -284 -2582 284 2582
<< labels >>
flabel metal1 11721 -7657 11721 -7657 0 FreeSans 400 0 0 0 vref_int
flabel metal1 27621 -7626 27621 -7626 0 FreeSans 400 0 0 0 vstart
flabel metal2 12874 -7070 12874 -7070 0 FreeSans 400 0 0 0 vbias_p
flabel metal2 12912 -7425 12912 -7425 0 FreeSans 400 0 0 0 vbias_c
flabel metal2 12820 -7931 12820 -7931 0 FreeSans 400 0 0 0 vbias_n
flabel metal3 10800 -6524 10800 -6524 0 FreeSans 400 0 0 0 vpass
flabel metal1 10194 -7632 10194 -7632 0 FreeSans 400 0 0 0 verr
flabel metal1 7903 -7803 7903 -7803 0 FreeSans 400 90 0 0 vm
flabel metal1 7447 -8672 7447 -8672 0 FreeSans 400 90 0 0 vref
flabel metal1 7346 -8991 7346 -8991 0 FreeSans 400 90 0 0 vref_int
flabel metal1 7039 -7713 7039 -7713 0 FreeSans 400 0 0 0 vx
flabel metal1 8350 -7725 8350 -7725 0 FreeSans 400 0 0 0 vy
flabel metal2 8258 -10049 8258 -10049 0 FreeSans 400 90 0 0 vref_ext
flabel metal2 27664 -6486 27664 -6486 0 FreeSans 400 0 0 0 vdd_start
flabel metal4 28188 -6478 28388 -6278 0 FreeSans 256 0 0 0 AVDD
port 0 nsew
flabel metal4 28225 -10398 28425 -10198 0 FreeSans 256 0 0 0 AVSS
port 2 nsew
flabel metal2 8176 -10750 8376 -10550 0 FreeSans 256 0 0 0 VREF_EXT
port 4 nsew
flabel metal2 9022 6637 9222 6837 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal2 8169 6695 8369 6895 0 FreeSans 256 0 0 0 SEL_EXT
port 5 nsew
flabel metal2 6055 6695 6255 6895 0 FreeSans 256 0 0 0 ENA
port 3 nsew
flabel metal2 8307 -9425 8307 -9425 0 FreeSans 400 0 0 0 nena
flabel metal1 6161 -8950 6161 -8950 0 FreeSans 400 90 0 0 sel_ext_3v3
flabel metal1 5737 -8932 5737 -8932 0 FreeSans 400 90 0 0 ena_3v3
flabel metal1 6744 -9430 6744 -9430 0 FreeSans 400 0 0 0 nsel_ext
<< end >>
